-------------------------------------------------------------------------------
--  HTLROM32                                                                 --
--  Copyright (C) 2002-2025 HT-LAB                                           --
--                                                                           --
-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- Project       :                                                           --
-- Purpose       :                                                           --
-- Library       :                                                           --
--                                                                           --
-- Created       : bin2text -vhd version  0.5                                --
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.ALL;

entity bootloader is
	port(clk    : in  std_logic;
		 abus   : in  std_logic_vector(12 downto 0);
		 ena    : in std_logic;
		 dbus   : out std_logic_vector(31 downto 0));
end bootloader;

architecture rtl of bootloader is
begin

	process(clk)
		begin
		if rising_edge(clk) then
			if ena='1' then
			case abus is
				when "0000000000000"  => dbus <= X"0001A801";
				when "0000000000001"  => dbus <= X"00000013";
				when "0000000000010"  => dbus <= X"00000013";
				when "0000000000011"  => dbus <= X"00000013";
				when "0000000000100"  => dbus <= X"00008137";
				when "0000000000101"  => dbus <= X"B8010113";
				when "0000000000110"  => dbus <= X"00002517";
				when "0000000000111"  => dbus <= X"15450513";
				when "0000000001000"  => dbus <= X"00000593";
				when "0000000001001"  => dbus <= X"01800613";
				when "0000000001010"  => dbus <= X"00C5D863";
				when "0000000001011"  => dbus <= X"C1944114";
				when "0000000001100"  => dbus <= X"05910511";
				when "0000000001101"  => dbus <= X"FEC5CCE3";
				when "0000000001110"  => dbus <= X"01800513";
				when "0000000001111"  => dbus <= X"02C00593";
				when "0000000010000"  => dbus <= X"00B55763";
				when "0000000010001"  => dbus <= X"00052023";
				when "0000000010010"  => dbus <= X"4DE30511";
				when "0000000010011"  => dbus <= X"10EFFEB5";
				when "0000000010100"  => dbus <= X"90024940";
				when "0000000010101"  => dbus <= X"00000000";
				when "0000000010110"  => dbus <= X"00000000";
				when "0000000010111"  => dbus <= X"00000000";
				when "0000000011000"  => dbus <= X"C04A1141";
				when "0000000011001"  => dbus <= X"01C52903";
				when "0000000011010"  => dbus <= X"C226C422";
				when "0000000011011"  => dbus <= X"842AC606";
				when "0000000011100"  => dbus <= X"02052C23";
				when "0000000011101"  => dbus <= X"02052E23";
				when "0000000011110"  => dbus <= X"99634481";
				when "0000000011111"  => dbus <= X"40B20124";
				when "0000000100000"  => dbus <= X"44924422";
				when "0000000100001"  => dbus <= X"45014902";
				when "0000000100010"  => dbus <= X"80820141";
				when "0000000100011"  => dbus <= X"85224585";
				when "0000000100100"  => dbus <= X"55832C55";
				when "0000000100101"  => dbus <= X"00EF0384";
				when "0000000100110"  => dbus <= X"1C233C10";
				when "0000000100111"  => dbus <= X"55FD02A4";
				when "0000000101000"  => dbus <= X"244D8522";
				when "0000000101001"  => dbus <= X"03845583";
				when "0000000101010"  => dbus <= X"3AF000EF";
				when "0000000101011"  => dbus <= X"02A41C23";
				when "0000000101100"  => dbus <= X"1D23E099";
				when "0000000101101"  => dbus <= X"048502A4";
				when "0000000101110"  => dbus <= X"E60DB7C9";
				when "0000000101111"  => dbus <= X"00051783";
				when "0000000110000"  => dbus <= X"F007F713";
				when "0000000110001"  => dbus <= X"83C107C2";
				when "0000000110010"  => dbus <= X"8FD983A1";
				when "0000000110011"  => dbus <= X"00F51023";
				when "0000000110100"  => dbus <= X"00059783";
				when "0000000110101"  => dbus <= X"F007F713";
				when "0000000110110"  => dbus <= X"83C107C2";
				when "0000000110111"  => dbus <= X"8FD983A1";
				when "0000000111000"  => dbus <= X"00F59023";
				when "0000000111001"  => dbus <= X"00251503";
				when "0000000111010"  => dbus <= X"00259783";
				when "0000000111011"  => dbus <= X"80828D1D";
				when "0000000111100"  => dbus <= X"CA261101";
				when "0000000111101"  => dbus <= X"00051483";
				when "0000000111110"  => dbus <= X"CC22CE06";
				when "0000000111111"  => dbus <= X"4074D793";
				when "0000001000000"  => dbus <= X"C64EC84A";
				when "0000001000001"  => dbus <= X"CB918B85";
				when "0000001000010"  => dbus <= X"07F4F513";
				when "0000001000011"  => dbus <= X"446240F2";
				when "0000001000100"  => dbus <= X"494244D2";
				when "0000001000101"  => dbus <= X"610549B2";
				when "0000001000110"  => dbus <= X"842E8082";
				when "0000001000111"  => dbus <= X"4034D593";
				when "0000001001000"  => dbus <= X"00F5F793";
				when "0000001001001"  => dbus <= X"00479593";
				when "0000001001010"  => dbus <= X"0074F713";
				when "0000001001011"  => dbus <= X"89AA8DDD";
				when "0000001001100"  => dbus <= X"03845783";
				when "0000001001101"  => dbus <= X"4685C31D";
				when "0000001001110"  => dbus <= X"1A638926";
				when "0000001001111"  => dbus <= X"863E04D7";
				when "0000001010000"  => dbus <= X"02840513";
				when "0000001010001"  => dbus <= X"57832F05";
				when "0000001010010"  => dbus <= X"191303C4";
				when "0000001010011"  => dbus <= X"59130105";
				when "0000001010100"  => dbus <= X"EF954109";
				when "0000001010101"  => dbus <= X"02A41E23";
				when "0000001010110"  => dbus <= X"0693A81D";
				when "0000001010111"  => dbus <= X"872E0220";
				when "0000001011000"  => dbus <= X"00D5D463";
				when "0000001011001"  => dbus <= X"02200713";
				when "0000001011010"  => dbus <= X"00241683";
				when "0000001011011"  => dbus <= X"00041603";
				when "0000001011100"  => dbus <= X"4C08484C";
				when "0000001011101"  => dbus <= X"0FF77713";
				when "0000001011110"  => dbus <= X"185000EF";
				when "0000001011111"  => dbus <= X"03E45783";
				when "0000001100000"  => dbus <= X"01051913";
				when "0000001100001"  => dbus <= X"41095913";
				when "0000001100010"  => dbus <= X"1F23E399";
				when "0000001100011"  => dbus <= X"558302A4";
				when "0000001100100"  => dbus <= X"15130384";
				when "0000001100101"  => dbus <= X"81410109";
				when "0000001100110"  => dbus <= X"2BF000EF";
				when "0000001100111"  => dbus <= X"02A41C23";
				when "0000001101000"  => dbus <= X"F004F493";
				when "0000001101001"  => dbus <= X"07F97513";
				when "0000001101010"  => dbus <= X"E4938CC9";
				when "0000001101011"  => dbus <= X"90230804";
				when "0000001101100"  => dbus <= X"BFA90099";
				when "0000001101101"  => dbus <= X"CA261101";
				when "0000001101110"  => dbus <= X"85B284AE";
				when "0000001101111"  => dbus <= X"CC22CE06";
				when "0000001110000"  => dbus <= X"373DC632";
				when "0000001110001"  => dbus <= X"842A4632";
				when "0000001110010"  => dbus <= X"85B28526";
				when "0000001110011"  => dbus <= X"05333715";
				when "0000001110100"  => dbus <= X"40F240A4";
				when "0000001110101"  => dbus <= X"44D24462";
				when "0000001110110"  => dbus <= X"80826105";
				when "0000001110111"  => dbus <= X"00059783";
				when "0000001111000"  => dbus <= X"00F51023";
				when "0000001111001"  => dbus <= X"00259783";
				when "0000001111010"  => dbus <= X"00F51123";
				when "0000001111011"  => dbus <= X"882A8082";
				when "0000001111100"  => dbus <= X"08934208";
				when "0000001111101"  => dbus <= X"FC630085";
				when "0000001111110"  => dbus <= X"429802E8";
				when "0000001111111"  => dbus <= X"00470313";
				when "0000010000000"  => dbus <= X"02F37763";
				when "0000010000001"  => dbus <= X"01162023";
				when "0000010000010"  => dbus <= X"00082783";
				when "0000010000011"  => dbus <= X"2023C11C";
				when "0000010000100"  => dbus <= X"C15800A8";
				when "0000010000101"  => dbus <= X"9703429C";
				when "0000010000110"  => dbus <= X"07910005";
				when "0000010000111"  => dbus <= X"415CC29C";
				when "0000010001000"  => dbus <= X"00E79023";
				when "0000010001001"  => dbus <= X"00259703";
				when "0000010001010"  => dbus <= X"00E79123";
				when "0000010001011"  => dbus <= X"45018082";
				when "0000010001100"  => dbus <= X"411C8082";
				when "0000010001101"  => dbus <= X"43D44158";
				when "0000010001110"  => dbus <= X"C3D8C154";
				when "0000010001111"  => dbus <= X"C1184398";
				when "0000010010000"  => dbus <= X"0007A023";
				when "0000010010001"  => dbus <= X"8082853E";
				when "0000010010010"  => dbus <= X"415841D4";
				when "0000010010011"  => dbus <= X"C1D8C154";
				when "0000010010100"  => dbus <= X"C1184198";
				when "0000010010101"  => dbus <= X"8082C188";
				when "0000010010110"  => dbus <= X"00259783";
				when "0000010010111"  => dbus <= X"0007DE63";
				when "0000010011000"  => dbus <= X"415CC115";
				when "0000010011001"  => dbus <= X"0007C703";
				when "0000010011010"  => dbus <= X"00059783";
				when "0000010011011"  => dbus <= X"00F71363";
				when "0000010011100"  => dbus <= X"41088082";
				when "0000010011101"  => dbus <= X"4108B7F5";
				when "0000010011110"  => dbus <= X"4158C511";
				when "0000010011111"  => dbus <= X"00271703";
				when "0000010100000"  => dbus <= X"FEF71BE3";
				when "0000010100001"  => dbus <= X"87AA8082";
				when "0000010100010"  => dbus <= X"E3914501";
				when "0000010100011"  => dbus <= X"43988082";
				when "0000010100100"  => dbus <= X"853EC388";
				when "0000010100101"  => dbus <= X"BFD587BA";
				when "0000010100110"  => dbus <= X"CC527179";
				when "0000010100111"  => dbus <= X"C462CA56";
				when "0000010101000"  => dbus <= X"C06AC266";
				when "0000010101001"  => dbus <= X"D422D606";
				when "0000010101010"  => dbus <= X"D04AD226";
				when "0000010101011"  => dbus <= X"C85ACE4E";
				when "0000010101100"  => dbus <= X"8C2EC65E";
				when "0000010101101"  => dbus <= X"8A2A8CB2";
				when "0000010101110"  => dbus <= X"4D054A85";
				when "0000010101111"  => dbus <= X"4B8184D2";
				when "0000010110000"  => dbus <= X"4A014B01";
				when "0000010110001"  => dbus <= X"2023E499";
				when "0000010110010"  => dbus <= X"5E63000B";
				when "0000010110011"  => dbus <= X"0A86057D";
				when "0000010110100"  => dbus <= X"0B85B7F5";
				when "0000010110101"  => dbus <= X"49018426";
				when "0000010110110"  => dbus <= X"09054000";
				when "0000010110111"  => dbus <= X"89D6E809";
				when "0000010111000"  => dbus <= X"00091A63";
				when "0000010111001"  => dbus <= X"00098363";
				when "0000010111010"  => dbus <= X"84A2E815";
				when "0000010111011"  => dbus <= X"95E3BFE1";
				when "0000010111100"  => dbus <= X"B7F5FF2A";
				when "0000010111101"  => dbus <= X"00098363";
				when "0000010111110"  => dbus <= X"87A2EC01";
				when "0000010111111"  => dbus <= X"40848426";
				when "0000011000000"  => dbus <= X"0063197D";
				when "0000011000001"  => dbus <= X"2023020B";
				when "0000011000010"  => dbus <= X"8B22008B";
				when "0000011000011"  => dbus <= X"BFC9843E";
				when "0000011000100"  => dbus <= X"40C8404C";
				when "0000011000101"  => dbus <= X"9C028666";
				when "0000011000110"  => dbus <= X"FEA051E3";
				when "0000011000111"  => dbus <= X"19FD401C";
				when "0000011001000"  => dbus <= X"8A22B7CD";
				when "0000011001001"  => dbus <= X"50B2B7DD";
				when "0000011001010"  => dbus <= X"85525422";
				when "0000011001011"  => dbus <= X"59025492";
				when "0000011001100"  => dbus <= X"4A6249F2";
				when "0000011001101"  => dbus <= X"4B424AD2";
				when "0000011001110"  => dbus <= X"4C224BB2";
				when "0000011001111"  => dbus <= X"4D024C92";
				when "0000011010000"  => dbus <= X"80826145";
				when "0000011010001"  => dbus <= X"C4A2715D";
				when "0000011010010"  => dbus <= X"5140D65E";
				when "0000011010011"  => dbus <= X"00451B83";
				when "0000011010100"  => dbus <= X"C0CAC2A6";
				when "0000011010101"  => dbus <= X"DA56DC52";
				when "0000011010110"  => dbus <= X"C686D85A";
				when "0000011010111"  => dbus <= X"862ADE4E";
				when "0000011011000"  => dbus <= X"1E238A2E";
				when "0000011011001"  => dbus <= X"1F230001";
				when "0000011011010"  => dbus <= X"4A8100B1";
				when "0000011011011"  => dbus <= X"49014B01";
				when "0000011011100"  => dbus <= X"CF634481";
				when "0000011011101"  => dbus <= X"090A077A";
				when "0000011011110"  => dbus <= X"41690933";
				when "0000011011111"  => dbus <= X"04C294CA";
				when "0000011100000"  => dbus <= X"596380C1";
				when "0000011100001"  => dbus <= X"05B70140";
				when "0000011100010"  => dbus <= X"85224000";
				when "0000011100011"  => dbus <= X"1B458593";
				when "0000011100100"  => dbus <= X"842A3721";
				when "0000011100101"  => dbus <= X"3D714008";
				when "0000011100110"  => dbus <= X"086C89AA";
				when "0000011100111"  => dbus <= X"3D6D8522";
				when "0000011101000"  => dbus <= X"E119892A";
				when "0000011101001"  => dbus <= X"00042903";
				when "0000011101010"  => dbus <= X"0C091763";
				when "0000011101011"  => dbus <= X"A703401C";
				when "0000011101100"  => dbus <= X"05B70049";
				when "0000011101101"  => dbus <= X"43D44000";
				when "0000011101110"  => dbus <= X"46018522";
				when "0000011101111"  => dbus <= X"00D9A223";
				when "0000011110000"  => dbus <= X"4398C3D8";
				when "0000011110001"  => dbus <= X"0BA58593";
				when "0000011110010"  => dbus <= X"00E9A023";
				when "0000011110011"  => dbus <= X"0137A023";
				when "0000011110100"  => dbus <= X"410035E1";
				when "0000011110101"  => dbus <= X"E855892A";
				when "0000011110110"  => dbus <= X"442640B6";
				when "0000011110111"  => dbus <= X"49068526";
				when "0000011111000"  => dbus <= X"59F24496";
				when "0000011111001"  => dbus <= X"5AD25A62";
				when "0000011111010"  => dbus <= X"5BB25B42";
				when "0000011111011"  => dbus <= X"80826161";
				when "0000011111100"  => dbus <= X"0FFAF793";
				when "0000011111101"  => dbus <= X"8522086C";
				when "0000011111110"  => dbus <= X"1E23C632";
				when "0000011111111"  => dbus <= X"3DA900F1";
				when "0000100000000"  => dbus <= X"852289AA";
				when "0000100000001"  => dbus <= X"842A3549";
				when "0000100000010"  => dbus <= X"9C634632";
				when "0000100000011"  => dbus <= X"411C0209";
				when "0000100000100"  => dbus <= X"0B420B05";
				when "0000100000101"  => dbus <= X"5B1343DC";
				when "0000100000110"  => dbus <= X"8783010B";
				when "0000100000111"  => dbus <= X"8B850017";
				when "0000100001000"  => dbus <= X"04C294BE";
				when "0000100001001"  => dbus <= X"178380C1";
				when "0000100001010"  => dbus <= X"C56301E1";
				when "0000100001011"  => dbus <= X"07850007";
				when "0000100001100"  => dbus <= X"00F11F23";
				when "0000100001101"  => dbus <= X"001A8793";
				when "0000100001110"  => dbus <= X"01079A93";
				when "0000100001111"  => dbus <= X"410ADA93";
				when "0000100010000"  => dbus <= X"A703BF0D";
				when "0000100010001"  => dbus <= X"09050049";
				when "0000100010010"  => dbus <= X"17830942";
				when "0000100010011"  => dbus <= X"59130007";
				when "0000100010100"  => dbus <= X"F7130109";
				when "0000100010101"  => dbus <= X"C7110017";
				when "0000100010110"  => dbus <= X"8B8587A5";
				when "0000100010111"  => dbus <= X"04C294BE";
				when "0000100011000"  => dbus <= X"A78380C1";
				when "0000100011001"  => dbus <= X"D3E10009";
				when "0000100011010"  => dbus <= X"A0234398";
				when "0000100011011"  => dbus <= X"401800E9";
				when "0000100011100"  => dbus <= X"C01CC398";
				when "0000100011101"  => dbus <= X"405CBF4D";
				when "0000100011110"  => dbus <= X"950385A6";
				when "0000100011111"  => dbus <= X"00EF0007";
				when "0000100100000"  => dbus <= X"84AA0110";
				when "0000100100001"  => dbus <= X"00092903";
				when "0000100100010"  => dbus <= X"2783B705";
				when "0000100100011"  => dbus <= X"85A60049";
				when "0000100100100"  => dbus <= X"00079503";
				when "0000100100101"  => dbus <= X"7FA000EF";
				when "0000100100110"  => dbus <= X"400084AA";
				when "0000100100111"  => dbus <= X"7139BF2D";
				when "0000100101000"  => dbus <= X"4451DC22";
				when "0000100101001"  => dbus <= X"02855433";
				when "0000100101010"  => dbus <= X"D84ADA26";
				when "0000100101011"  => dbus <= X"D452D64E";
				when "0000100101100"  => dbus <= X"DE06D256";
				when "0000100101101"  => dbus <= X"A02377E1";
				when "0000100101110"  => dbus <= X"87930005";
				when "0000100101111"  => dbus <= X"89AE0807";
				when "0000100110000"  => dbus <= X"08348932";
				when "0000100110001"  => dbus <= X"854E0070";
				when "0000100110010"  => dbus <= X"14794A01";
				when "0000100110011"  => dbus <= X"00341493";
				when "0000100110100"  => dbus <= X"C1C494AE";
				when "0000100110101"  => dbus <= X"00F49023";
				when "0000100110110"  => dbus <= X"00049123";
				when "0000100110111"  => dbus <= X"00858793";
				when "0000100111000"  => dbus <= X"8793C63E";
				when "0000100111001"  => dbus <= X"CC3E0044";
				when "0000100111010"  => dbus <= X"00241A93";
				when "0000100111011"  => dbus <= X"800007B7";
				when "0000100111100"  => dbus <= X"FFF7C793";
				when "0000100111101"  => dbus <= X"CE3E9AA6";
				when "0000100111110"  => dbus <= X"87D68726";
				when "0000100111111"  => dbus <= X"39C5086C";
				when "0000101000000"  => dbus <= X"028A6C63";
				when "0000101000001"  => dbus <= X"54334515";
				when "0000101000010"  => dbus <= X"A78302A4";
				when "0000101000011"  => dbus <= X"66110009";
				when "0000101000100"  => dbus <= X"167D4705";
				when "0000101000101"  => dbus <= X"E9A9438C";
				when "0000101000110"  => dbus <= X"400005B7";
				when "0000101000111"  => dbus <= X"4601854E";
				when "0000101001000"  => dbus <= X"0BA58593";
				when "0000101001001"  => dbus <= X"50F23B95";
				when "0000101001010"  => dbus <= X"54D25462";
				when "0000101001011"  => dbus <= X"59B25942";
				when "0000101001100"  => dbus <= X"5A925A22";
				when "0000101001101"  => dbus <= X"80826121";
				when "0000101001110"  => dbus <= X"010A1713";
				when "0000101001111"  => dbus <= X"47B38341";
				when "0000101010000"  => dbus <= X"078E0127";
				when "0000101010001"  => dbus <= X"F7938B1D";
				when "0000101010010"  => dbus <= X"8FD90787";
				when "0000101010011"  => dbus <= X"00879713";
				when "0000101010100"  => dbus <= X"1E238FD9";
				when "0000101010101"  => dbus <= X"872600F1";
				when "0000101010110"  => dbus <= X"083487D6";
				when "0000101010111"  => dbus <= X"086C0070";
				when "0000101011000"  => dbus <= X"3171854E";
				when "0000101011001"  => dbus <= X"BF690A05";
				when "0000101011010"  => dbus <= X"776343C8";
				when "0000101011011"  => dbus <= X"11230087";
				when "0000101011100"  => dbus <= X"070500E5";
				when "0000101011101"  => dbus <= X"BF7987AE";
				when "0000101011110"  => dbus <= X"01071693";
				when "0000101011111"  => dbus <= X"879382C1";
				when "0000101100000"  => dbus <= X"07A20016";
				when "0000101100001"  => dbus <= X"7007F793";
				when "0000101100010"  => dbus <= X"0126C6B3";
				when "0000101100011"  => dbus <= X"8FF18FD5";
				when "0000101100100"  => dbus <= X"00F51123";
				when "0000101100101"  => dbus <= X"1141BFF9";
				when "0000101100110"  => dbus <= X"E211C622";
				when "0000101100111"  => dbus <= X"47014605";
				when "0000101101000"  => dbus <= X"A0294781";
				when "0000101101001"  => dbus <= X"87330785";
				when "0000101101010"  => dbus <= X"070E02F7";
				when "0000101101011"  => dbus <= X"FEA76CE3";
				when "0000101101100"  => dbus <= X"FFF78513";
				when "0000101101101"  => dbus <= X"02A507B3";
				when "0000101101110"  => dbus <= X"99F115FD";
				when "0000101101111"  => dbus <= X"12930591";
				when "0000101110000"  => dbus <= X"4E810015";
				when "0000101110001"  => dbus <= X"63C14F05";
				when "0000101110010"  => dbus <= X"00179893";
				when "0000101110011"  => dbus <= X"011587B3";
				when "0000101110100"  => dbus <= X"84338FBE";
				when "0000101110101"  => dbus <= X"EC6340F5";
				when "0000101110110"  => dbus <= X"C69C04AE";
				when "0000101110111"  => dbus <= X"17FD97C6";
				when "0000101111000"  => dbus <= X"9BF14432";
				when "0000101111001"  => dbus <= X"C2CC0791";
				when "0000101111010"  => dbus <= X"C288C6DC";
				when "0000101111011"  => dbus <= X"80820141";
				when "0000101111100"  => dbus <= X"02E60633";
				when "0000101111101"  => dbus <= X"01071813";
				when "0000101111110"  => dbus <= X"01085813";
				when "0000101111111"  => dbus <= X"66330305";
				when "0000110000000"  => dbus <= X"07330276";
				when "0000110000001"  => dbus <= X"074200C8";
				when "0000110000010"  => dbus <= X"10238341";
				when "0000110000011"  => dbus <= X"974200EE";
				when "0000110000100"  => dbus <= X"0FF77713";
				when "0000110000101"  => dbus <= X"01C40833";
				when "0000110000110"  => dbus <= X"00E81023";
				when "0000110000111"  => dbus <= X"07330E09";
				when "0000110001000"  => dbus <= X"67E301E3";
				when "0000110001001"  => dbus <= X"0E85FCA3";
				when "0000110001010"  => dbus <= X"9F2A9F96";
				when "0000110001011"  => dbus <= X"8E7EB76D";
				when "0000110001100"  => dbus <= X"B7F54301";
				when "0000110001101"  => dbus <= X"00251E93";
				when "0000110001110"  => dbus <= X"47814801";
				when "0000110001111"  => dbus <= X"47014681";
				when "0000110010000"  => dbus <= X"02A81D63";
				when "0000110010001"  => dbus <= X"8082853E";
				when "0000110010010"  => dbus <= X"00032E03";
				when "0000110010011"  => dbus <= X"83C107C2";
				when "0000110010100"  => dbus <= X"5E639772";
				when "0000110010101"  => dbus <= X"07A900E6";
				when "0000110010110"  => dbus <= X"87C107C2";
				when "0000110010111"  => dbus <= X"08854701";
				when "0000110011000"  => dbus <= X"86F20311";
				when "0000110011001"  => dbus <= X"FEA892E3";
				when "0000110011010"  => dbus <= X"95F60805";
				when "0000110011011"  => dbus <= X"A6B3BFD1";
				when "0000110011100"  => dbus <= X"97B601C6";
				when "0000110011101"  => dbus <= X"87C107C2";
				when "0000110011110"  => dbus <= X"832EB7DD";
				when "0000110011111"  => dbus <= X"B7DD4881";
				when "0000110100000"  => dbus <= X"00151E13";
				when "0000110100001"  => dbus <= X"00251E93";
				when "0000110100010"  => dbus <= X"92634781";
				when "0000110100011"  => dbus <= X"808202A7";
				when "0000110100100"  => dbus <= X"00081303";
				when "0000110100101"  => dbus <= X"08090705";
				when "0000110100110"  => dbus <= X"02D30333";
				when "0000110100111"  => dbus <= X"AE230891";
				when "0000110101000"  => dbus <= X"17E3FE68";
				when "0000110101001"  => dbus <= X"0785FEA7";
				when "0000110101010"  => dbus <= X"95F69672";
				when "0000110101011"  => dbus <= X"88AEBFF9";
				when "0000110101100"  => dbus <= X"47018832";
				when "0000110101101"  => dbus <= X"1893B7FD";
				when "0000110101110"  => dbus <= X"47010015";
				when "0000110101111"  => dbus <= X"00A71F63";
				when "0000110110000"  => dbus <= X"D8038082";
				when "0000110110001"  => dbus <= X"06850007";
				when "0000110110010"  => dbus <= X"98320789";
				when "0000110110011"  => dbus <= X"FF079F23";
				when "0000110110100"  => dbus <= X"FEA699E3";
				when "0000110110101"  => dbus <= X"95C60705";
				when "0000110110110"  => dbus <= X"87AEB7D5";
				when "0000110110111"  => dbus <= X"BFCD4681";
				when "0000110111000"  => dbus <= X"00151893";
				when "0000110111001"  => dbus <= X"952E050A";
				when "0000110111010"  => dbus <= X"00B51363";
				when "0000110111011"  => dbus <= X"47818082";
				when "0000110111100"  => dbus <= X"08334701";
				when "0000110111101"  => dbus <= X"833300F6";
				when "0000110111110"  => dbus <= X"180300F6";
				when "0000110111111"  => dbus <= X"13030008";
				when "0000111000000"  => dbus <= X"07890003";
				when "0000111000001"  => dbus <= X"02680833";
				when "0000111000010"  => dbus <= X"94E39742";
				when "0000111000011"  => dbus <= X"C198FEF8";
				when "0000111000100"  => dbus <= X"05919646";
				when "0000111000101"  => dbus <= X"1293BFD1";
				when "0000111000110"  => dbus <= X"1F930025";
				when "0000111000111"  => dbus <= X"48010015";
				when "0000111001000"  => dbus <= X"02A81F63";
				when "0000111001001"  => dbus <= X"17938082";
				when "0000111001010"  => dbus <= X"97B60017";
				when "0000111001011"  => dbus <= X"43018EB2";
				when "0000111001100"  => dbus <= X"9F034E01";
				when "0000111001101"  => dbus <= X"9383000E";
				when "0000111001110"  => dbus <= X"0E050007";
				when "0000111001111"  => dbus <= X"0F330E89";
				when "0000111010000"  => dbus <= X"97FE027F";
				when "0000111010001"  => dbus <= X"16E3937A";
				when "0000111010010"  => dbus <= X"A023FFC5";
				when "0000111010011"  => dbus <= X"07050068";
				when "0000111010100"  => dbus <= X"1AE30891";
				when "0000111010101"  => dbus <= X"0805FCA7";
				when "0000111010110"  => dbus <= X"967E9596";
				when "0000111010111"  => dbus <= X"88AEB7D1";
				when "0000111011000"  => dbus <= X"BFC54701";
				when "0000111011001"  => dbus <= X"00251393";
				when "0000111011010"  => dbus <= X"00151293";
				when "0000111011011"  => dbus <= X"18634301";
				when "0000111011100"  => dbus <= X"808204A3";
				when "0000111011101"  => dbus <= X"00189713";
				when "0000111011110"  => dbus <= X"8FB29736";
				when "0000111011111"  => dbus <= X"4F014E81";
				when "0000111100000"  => dbus <= X"00071803";
				when "0000111100001"  => dbus <= X"000F9783";
				when "0000111100010"  => dbus <= X"0F890F05";
				when "0000111100011"  => dbus <= X"030787B3";
				when "0000111100100"  => dbus <= X"D8139716";
				when "0000111100101"  => dbus <= X"87954027";
				when "0000111100110"  => dbus <= X"00F87813";
				when "0000111100111"  => dbus <= X"07F7F793";
				when "0000111101000"  => dbus <= X"02F807B3";
				when "0000111101001"  => dbus <= X"1DE39EBE";
				when "0000111101010"  => dbus <= X"2023FDE5";
				when "0000111101011"  => dbus <= X"088501DE";
				when "0000111101100"  => dbus <= X"91E30E11";
				when "0000111101101"  => dbus <= X"0305FCA8";
				when "0000111101110"  => dbus <= X"9616959E";
				when "0000111101111"  => dbus <= X"8E2EBF4D";
				when "0000111110000"  => dbus <= X"BFC54881";
				when "0000111110001"  => dbus <= X"C84A1101";
				when "0000111110010"  => dbus <= X"CA268932";
				when "0000111110011"  => dbus <= X"C452863A";
				when "0000111110100"  => dbus <= X"7A7D84AE";
				when "0000111110101"  => dbus <= X"CE0685CA";
				when "0000111110110"  => dbus <= X"01476A33";
				when "0000111110111"  => dbus <= X"C64ECC22";
				when "0000111111000"  => dbus <= X"89BAC256";
				when "0000111111001"  => dbus <= X"842AC05A";
				when "0000111111010"  => dbus <= X"35F18AB6";
				when "0000111111011"  => dbus <= X"864A86CE";
				when "0000111111100"  => dbus <= X"852285A6";
				when "0000111111101"  => dbus <= X"86523571";
				when "0000111111110"  => dbus <= X"852285A6";
				when "0000111111111"  => dbus <= X"45813D25";
				when "0001000000000"  => dbus <= X"86D62179";
				when "0001000000001"  => dbus <= X"864A8B2A";
				when "0001000000010"  => dbus <= X"852285A6";
				when "0001000000011"  => dbus <= X"86523DD1";
				when "0001000000100"  => dbus <= X"852285A6";
				when "0001000000101"  => dbus <= X"85DA3505";
				when "0001000000110"  => dbus <= X"86D6299D";
				when "0001000000111"  => dbus <= X"864A8B2A";
				when "0001000001000"  => dbus <= X"852285A6";
				when "0001000001001"  => dbus <= X"86523DCD";
				when "0001000001010"  => dbus <= X"852285A6";
				when "0001000001011"  => dbus <= X"85DA3521";
				when "0001000001100"  => dbus <= X"86D629B9";
				when "0001000001101"  => dbus <= X"864A8B2A";
				when "0001000001110"  => dbus <= X"852285A6";
				when "0001000001111"  => dbus <= X"86523725";
				when "0001000010000"  => dbus <= X"852285A6";
				when "0001000010001"  => dbus <= X"85DA3BC5";
				when "0001000010010"  => dbus <= X"06332199";
				when "0001000010011"  => dbus <= X"06424130";
				when "0001000010100"  => dbus <= X"85CA84AA";
				when "0001000010101"  => dbus <= X"86418522";
				when "0001000010110"  => dbus <= X"40F23DB9";
				when "0001000010111"  => dbus <= X"95134462";
				when "0001000011000"  => dbus <= X"49420104";
				when "0001000011001"  => dbus <= X"49B244D2";
				when "0001000011010"  => dbus <= X"4A924A22";
				when "0001000011011"  => dbus <= X"85414B02";
				when "0001000011100"  => dbus <= X"80826105";
				when "0001000011101"  => dbus <= X"C4221141";
				when "0001000011110"  => dbus <= X"8432872E";
				when "0001000011111"  => dbus <= X"4514454C";
				when "0001000100000"  => dbus <= X"41084150";
				when "0001000100001"  => dbus <= X"3F3DC606";
				when "0001000100010"  => dbus <= X"442285A2";
				when "0001000100011"  => dbus <= X"014140B2";
				when "0001000100100"  => dbus <= X"1141AEFD";
				when "0001000100101"  => dbus <= X"00EFC606";
				when "0001000100110"  => dbus <= X"40B22F10";
				when "0001000100111"  => dbus <= X"812105E2";
				when "0001000101000"  => dbus <= X"01418D4D";
				when "0001000101001"  => dbus <= X"11418082";
				when "0001000101010"  => dbus <= X"37E5C606";
				when "0001000101011"  => dbus <= X"2E2340B2";
				when "0001000101100"  => dbus <= X"85AA00A0";
				when "0001000101101"  => dbus <= X"40002537";
				when "0001000101110"  => dbus <= X"01450513";
				when "0001000101111"  => dbus <= X"AB510141";
				when "0001000110000"  => dbus <= X"C6061141";
				when "0001000110001"  => dbus <= X"40B237F9";
				when "0001000110010"  => dbus <= X"00A02C23";
				when "0001000110011"  => dbus <= X"253785AA";
				when "0001000110100"  => dbus <= X"05134000";
				when "0001000110101"  => dbus <= X"01410245";
				when "0001000110110"  => dbus <= X"2503ABAD";
				when "0001000110111"  => dbus <= X"27830180";
				when "0001000111000"  => dbus <= X"8D1D01C0";
				when "0001000111001"  => dbus <= X"07938082";
				when "0001000111010"  => dbus <= X"55330B70";
				when "0001000111011"  => dbus <= X"808202F5";
				when "0001000111100"  => dbus <= X"C4221141";
				when "0001000111101"  => dbus <= X"2537842A";
				when "0001000111110"  => dbus <= X"05134000";
				when "0001000111111"  => dbus <= X"C6060345";
				when "0001001000000"  => dbus <= X"47852B89";
				when "0001001000001"  => dbus <= X"00F40023";
				when "0001001000010"  => dbus <= X"442240B2";
				when "0001001000011"  => dbus <= X"80820141";
				when "0001001000100"  => dbus <= X"00050023";
				when "0001001000101"  => dbus <= X"47818082";
				when "0001001000110"  => dbus <= X"05854681";
				when "0001001000111"  => dbus <= X"00F68333";
				when "0001001001000"  => dbus <= X"283705C2";
				when "0001001001001"  => dbus <= X"2E374000";
				when "0001001001010"  => dbus <= X"0F134000";
				when "0001001001011"  => dbus <= X"0393FFF5";
				when "0001001001100"  => dbus <= X"81C10013";
				when "0001001001101"  => dbus <= X"0F934701";
				when "0001001001110"  => dbus <= X"429102C0";
				when "0001001001111"  => dbus <= X"BA080813";
				when "0001001010000"  => dbus <= X"B6CE0E13";
				when "0001001010001"  => dbus <= X"05E3E963";
				when "0001001010010"  => dbus <= X"04A6E163";
				when "0001001010011"  => dbus <= X"97C28082";
				when "0001001010100"  => dbus <= X"47914398";
				when "0001001010101"  => dbus <= X"83330585";
				when "0001001010110"  => dbus <= X"05C200F6";
				when "0001001010111"  => dbus <= X"00130393";
				when "0001001011000"  => dbus <= X"EC6381C1";
				when "0001001011001"  => dbus <= X"EC6303E3";
				when "0001001011010"  => dbus <= X"443200A6";
				when "0001001011011"  => dbus <= X"80820141";
				when "0001001011100"  => dbus <= X"47A14B98";
				when "0001001011101"  => dbus <= X"5398B7C5";
				when "0001001011110"  => dbus <= X"5B98BFED";
				when "0001001011111"  => dbus <= X"07B3BFDD";
				when "0001001100000"  => dbus <= X"802300D6";
				when "0001001100001"  => dbus <= X"06850007";
				when "0001001100010"  => dbus <= X"07B3BFF9";
				when "0001001100011"  => dbus <= X"802300D6";
				when "0001001100100"  => dbus <= X"06850007";
				when "0001001100101"  => dbus <= X"1141BF55";
				when "0001001100110"  => dbus <= X"C395C622";
				when "0001001100111"  => dbus <= X"0EB34881";
				when "0001001101000"  => dbus <= X"C4030117";
				when "0001001101001"  => dbus <= X"8EB3000E";
				when "0001001101010"  => dbus <= X"9EB20116";
				when "0001001101011"  => dbus <= X"008E8023";
				when "0001001101100"  => dbus <= X"96E30885";
				when "0001001101101"  => dbus <= X"9332FF17";
				when "0001001101110"  => dbus <= X"01F30023";
				when "0001001101111"  => dbus <= X"F713869E";
				when "0001001110000"  => dbus <= X"17750075";
				when "0001001110001"  => dbus <= X"D7930742";
				when "0001001110010"  => dbus <= X"83410015";
				when "0001001110011"  => dbus <= X"E0E38BB1";
				when "0001001110100"  => dbus <= X"070AF8E2";
				when "0001001110101"  => dbus <= X"43189772";
				when "0001001110110"  => dbus <= X"870297C2";
				when "0001001110111"  => dbus <= X"28374114";
				when "0001001111000"  => dbus <= X"47014000";
				when "0001001111001"  => dbus <= X"0E134305";
				when "0001001111010"  => dbus <= X"4E9D02C0";
				when "0001001111011"  => dbus <= X"B8080813";
				when "0001001111100"  => dbus <= X"0F134625";
				when "0001001111101"  => dbus <= X"08930450";
				when "0001001111110"  => dbus <= X"C78302E0";
				when "0001001111111"  => dbus <= X"C3990006";
				when "0001010000000"  => dbus <= X"00671563";
				when "0001010000001"  => dbus <= X"853AC114";
				when "0001010000010"  => dbus <= X"06858082";
				when "0001010000011"  => dbus <= X"FFC78CE3";
				when "0001010000100"  => dbus <= X"FEEEE5E3";
				when "0001010000101"  => dbus <= X"00271F93";
				when "0001010000110"  => dbus <= X"AF839FC2";
				when "0001010000111"  => dbus <= X"8F82000F";
				when "0001010001000"  => dbus <= X"FD078F93";
				when "0001010001001"  => dbus <= X"0FFFFF93";
				when "0001010001010"  => dbus <= X"70634711";
				when "0001010001011"  => dbus <= X"8F9303F6";
				when "0001010001100"  => dbus <= X"FF93FD57";
				when "0001010001101"  => dbus <= X"47090FDF";
				when "0001010001110"  => dbus <= X"000F8963";
				when "0001010001111"  => dbus <= X"86634715";
				when "0001010010000"  => dbus <= X"41DC0117";
				when "0001010010001"  => dbus <= X"07854705";
				when "0001010010010"  => dbus <= X"419CC1DC";
				when "0001010010011"  => dbus <= X"C19C0785";
				when "0001010010100"  => dbus <= X"4598B76D";
				when "0001010010101"  => dbus <= X"FD078F93";
				when "0001010010110"  => dbus <= X"0FFFFF93";
				when "0001010010111"  => dbus <= X"77630705";
				when "0001010011000"  => dbus <= X"986301F6";
				when "0001010011001"  => dbus <= X"C5980117";
				when "0001010011010"  => dbus <= X"BF414715";
				when "0001010011011"  => dbus <= X"4711C598";
				when "0001010011100"  => dbus <= X"C598B769";
				when "0001010011101"  => dbus <= X"B7514705";
				when "0001010011110"  => dbus <= X"01179663";
				when "0001010011111"  => dbus <= X"0785499C";
				when "0001010100000"  => dbus <= X"B7DDC99C";
				when "0001010100001"  => dbus <= X"FD078793";
				when "0001010100010"  => dbus <= X"0FF7F793";
				when "0001010100011"  => dbus <= X"F6F677E3";
				when "0001010100100"  => dbus <= X"0785499C";
				when "0001010100101"  => dbus <= X"BFF9C99C";
				when "0001010100110"  => dbus <= X"0DF7FF93";
				when "0001010100111"  => dbus <= X"01EF9763";
				when "0001010101000"  => dbus <= X"470D49DC";
				when "0001010101001"  => dbus <= X"C9DC0785";
				when "0001010101010"  => dbus <= X"8793BF89";
				when "0001010101011"  => dbus <= X"F793FD07";
				when "0001010101100"  => dbus <= X"74E30FF7";
				when "0001010101101"  => dbus <= X"49DCF4F6";
				when "0001010101110"  => dbus <= X"C9DC0785";
				when "0001010101111"  => dbus <= X"45D8BF65";
				when "0001010110000"  => dbus <= X"FD578793";
				when "0001010110001"  => dbus <= X"0FD7F793";
				when "0001010110010"  => dbus <= X"C5D80705";
				when "0001010110011"  => dbus <= X"F3DD4719";
				when "0001010110100"  => dbus <= X"4D98B72D";
				when "0001010110101"  => dbus <= X"FD078793";
				when "0001010110110"  => dbus <= X"0FF7F793";
				when "0001010110111"  => dbus <= X"CD980705";
				when "0001010111000"  => dbus <= X"7CE3471D";
				when "0001010111001"  => dbus <= X"B779F0F6";
				when "0001010111010"  => dbus <= X"FD078793";
				when "0001010111011"  => dbus <= X"0FF7F793";
				when "0001010111100"  => dbus <= X"F0F675E3";
				when "0001010111101"  => dbus <= X"078541DC";
				when "0001010111110"  => dbus <= X"BFADC1DC";
				when "0001010111111"  => dbus <= X"DCA27119";
				when "0001011000000"  => dbus <= X"D8CADAA6";
				when "0001011000001"  => dbus <= X"D4D2D6CE";
				when "0001011000010"  => dbus <= X"893E842E";
				when "0001011000011"  => dbus <= X"DE86CE2E";
				when "0001011000100"  => dbus <= X"8A3684AA";
				when "0001011000101"  => dbus <= X"458189BA";
				when "0001011000110"  => dbus <= X"02000793";
				when "0001011000111"  => dbus <= X"972E0098";
				when "0001011001000"  => dbus <= X"00072023";
				when "0001011001001"  => dbus <= X"972E1018";
				when "0001011001010"  => dbus <= X"00072023";
				when "0001011001011"  => dbus <= X"97E30591";
				when "0001011001100"  => dbus <= X"47F2FEF5";
				when "0001011001101"  => dbus <= X"0007C783";
				when "0001011001110"  => dbus <= X"CE22EFA1";
				when "0001011001111"  => dbus <= X"071394A2";
				when "0001011010000"  => dbus <= X"47F202C0";
				when "0001011010001"  => dbus <= X"0697E463";
				when "0001011010010"  => dbus <= X"47F2CE22";
				when "0001011010011"  => dbus <= X"0007C783";
				when "0001011010100"  => dbus <= X"CE22EBAD";
				when "0001011010101"  => dbus <= X"02C00713";
				when "0001011010110"  => dbus <= X"E06347F2";
				when "0001011010111"  => dbus <= X"44010897";
				when "0001011011000"  => dbus <= X"02000493";
				when "0001011011001"  => dbus <= X"97A2101C";
				when "0001011011010"  => dbus <= X"85CA4388";
				when "0001011011011"  => dbus <= X"009C2219";
				when "0001011011100"  => dbus <= X"85AA97A2";
				when "0001011011101"  => dbus <= X"04114388";
				when "0001011011110"  => dbus <= X"892A28ED";
				when "0001011011111"  => dbus <= X"FE9414E3";
				when "0001011100000"  => dbus <= X"546650F6";
				when "0001011100001"  => dbus <= X"594654D6";
				when "0001011100010"  => dbus <= X"5A2659B6";
				when "0001011100011"  => dbus <= X"80826109";
				when "0001011100100"  => dbus <= X"0868008C";
				when "0001011100101"  => dbus <= X"3599C632";
				when "0001011100110"  => dbus <= X"050A109C";
				when "0001011100111"  => dbus <= X"2783953E";
				when "0001011101000"  => dbus <= X"4632FC05";
				when "0001011101001"  => dbus <= X"20230785";
				when "0001011101010"  => dbus <= X"B761FCF5";
				when "0001011101011"  => dbus <= X"0007C583";
				when "0001011101100"  => dbus <= X"00E58563";
				when "0001011101101"  => dbus <= X"80238DB1";
				when "0001011101110"  => dbus <= X"47F200B7";
				when "0001011101111"  => dbus <= X"CE3E97CE";
				when "0001011110000"  => dbus <= X"008CB749";
				when "0001011110001"  => dbus <= X"3D190868";
				when "0001011110010"  => dbus <= X"050A109C";
				when "0001011110011"  => dbus <= X"2783953E";
				when "0001011110100"  => dbus <= X"0785FC05";
				when "0001011110101"  => dbus <= X"FCF52023";
				when "0001011110110"  => dbus <= X"C603BF8D";
				when "0001011110111"  => dbus <= X"06630007";
				when "0001011111000"  => dbus <= X"463300E6";
				when "0001011111001"  => dbus <= X"80230146";
				when "0001011111010"  => dbus <= X"47F200C7";
				when "0001011111011"  => dbus <= X"CE3E97CE";
				when "0001011111100"  => dbus <= X"157DB7A5";
				when "0001011111101"  => dbus <= X"E9634791";
				when "0001011111110"  => dbus <= X"27B702A7";
				when "0001011111111"  => dbus <= X"87934000";
				when "0001100000000"  => dbus <= X"050ABE07";
				when "0001100000001"  => dbus <= X"411C953E";
				when "0001100000010"  => dbus <= X"25038782";
				when "0001100000011"  => dbus <= X"80820280";
				when "0001100000100"  => dbus <= X"02402503";
				when "0001100000101"  => dbus <= X"25038082";
				when "0001100000110"  => dbus <= X"80820140";
				when "0001100000111"  => dbus <= X"01002503";
				when "0001100001000"  => dbus <= X"25038082";
				when "0001100001001"  => dbus <= X"80820200";
				when "0001100001010"  => dbus <= X"80824501";
				when "0001100001011"  => dbus <= X"47A16691";
				when "0001100001100"  => dbus <= X"76610689";
				when "0001100001101"  => dbus <= X"00A5C733";
				when "0001100001110"  => dbus <= X"81058B05";
				when "0001100001111"  => dbus <= X"8DB5C311";
				when "0001100010000"  => dbus <= X"C7018185";
				when "0001100010001"  => dbus <= X"05C28DD1";
				when "0001100010010"  => dbus <= X"17FD81C1";
				when "0001100010011"  => dbus <= X"0FF7F793";
				when "0001100010100"  => dbus <= X"852EF3F5";
				when "0001100010101"  => dbus <= X"11418082";
				when "0001100010110"  => dbus <= X"842AC422";
				when "0001100010111"  => dbus <= X"0FF57513";
				when "0001100011000"  => dbus <= X"37E9C606";
				when "0001100011001"  => dbus <= X"551385AA";
				when "0001100011010"  => dbus <= X"44220084";
				when "0001100011011"  => dbus <= X"014140B2";
				when "0001100011100"  => dbus <= X"1141BF75";
				when "0001100011101"  => dbus <= X"842AC422";
				when "0001100011110"  => dbus <= X"81410542";
				when "0001100011111"  => dbus <= X"3FE1C606";
				when "0001100100000"  => dbus <= X"551385AA";
				when "0001100100001"  => dbus <= X"44220104";
				when "0001100100010"  => dbus <= X"014140B2";
				when "0001100100011"  => dbus <= X"0542B7E9";
				when "0001100100100"  => dbus <= X"B7D18141";
				when "0001100100101"  => dbus <= X"80824501";
				when "0001100100110"  => dbus <= X"0407F813";
				when "0001100100111"  => dbus <= X"0E63715D";
				when "0001100101000"  => dbus <= X"28B70008";
				when "0001100101001"  => dbus <= X"88934000";
				when "0001100101010"  => dbus <= X"FF931288";
				when "0001100101011"  => dbus <= X"8B630107";
				when "0001100101100"  => dbus <= X"9BF9000F";
				when "0001100101101"  => dbus <= X"02000E13";
				when "0001100101110"  => dbus <= X"28B7A821";
				when "0001100101111"  => dbus <= X"88934000";
				when "0001100110000"  => dbus <= X"B7E51008";
				when "0001100110001"  => dbus <= X"0017F813";
				when "0001100110010"  => dbus <= X"03000E13";
				when "0001100110011"  => dbus <= X"FE0804E3";
				when "0001100110100"  => dbus <= X"0027F813";
				when "0001100110101"  => dbus <= X"09634301";
				when "0001100110110"  => dbus <= X"D1630008";
				when "0001100110111"  => dbus <= X"05B30605";
				when "0001100111000"  => dbus <= X"16FD40B0";
				when "0001100111001"  => dbus <= X"02D00313";
				when "0001100111010"  => dbus <= X"0207F293";
				when "0001100111011"  => dbus <= X"00028663";
				when "0001100111100"  => dbus <= X"15634841";
				when "0001100111101"  => dbus <= X"16F90706";
				when "0001100111110"  => dbus <= X"0593E5BD";
				when "0001100111111"  => dbus <= X"06230300";
				when "0001101000000"  => dbus <= X"480500B1";
				when "0001101000001"  => dbus <= X"536385C2";
				when "0001101000010"  => dbus <= X"85BA00E8";
				when "0001101000011"  => dbus <= X"8E8D8BC5";
				when "0001101000100"  => dbus <= X"0563CFC1";
				when "0001101000101"  => dbus <= X"00230003";
				when "0001101000110"  => dbus <= X"05050065";
				when "0001101000111"  => dbus <= X"00028A63";
				when "0001101001000"  => dbus <= X"196347A1";
				when "0001101001001"  => dbus <= X"079308F6";
				when "0001101001010"  => dbus <= X"00230300";
				when "0001101001011"  => dbus <= X"050500F5";
				when "0001101001100"  => dbus <= X"0A0F8E63";
				when "0001101001101"  => dbus <= X"071395AA";
				when "0001101001110"  => dbus <= X"A0C10300";
				when "0001101001111"  => dbus <= X"0047F813";
				when "0001101010000"  => dbus <= X"00080663";
				when "0001101010001"  => dbus <= X"031316FD";
				when "0001101010010"  => dbus <= X"BF7902B0";
				when "0001101010011"  => dbus <= X"0087F813";
				when "0001101010100"  => dbus <= X"F8080CE3";
				when "0001101010101"  => dbus <= X"031316FD";
				when "0001101010110"  => dbus <= X"B7790200";
				when "0001101010111"  => dbus <= X"1DE34821";
				when "0001101011000"  => dbus <= X"16FDF906";
				when "0001101011001"  => dbus <= X"0E93BF51";
				when "0001101011010"  => dbus <= X"480100C1";
				when "0001101011011"  => dbus <= X"02C5FF33";
				when "0001101011100"  => dbus <= X"080583AE";
				when "0001101011101"  => dbus <= X"9F460E85";
				when "0001101011110"  => dbus <= X"000F4F03";
				when "0001101011111"  => dbus <= X"02C5D5B3";
				when "0001101100000"  => dbus <= X"FFEE8FA3";
				when "0001101100001"  => dbus <= X"FEC3F4E3";
				when "0001101100010"  => dbus <= X"0785BFB5";
				when "0001101100011"  => dbus <= X"FFD78FA3";
				when "0001101100100"  => dbus <= X"40F88733";
				when "0001101100101"  => dbus <= X"FEE04BE3";
				when "0001101100110"  => dbus <= X"D36387B6";
				when "0001101100111"  => dbus <= X"47810006";
				when "0001101101000"  => dbus <= X"953E16FD";
				when "0001101101001"  => dbus <= X"B7B58E9D";
				when "0001101101010"  => dbus <= X"08B387AA";
				when "0001101101011"  => dbus <= X"0E9300D5";
				when "0001101101100"  => dbus <= X"BFF90200";
				when "0001101101101"  => dbus <= X"1DE347C1";
				when "0001101101110"  => dbus <= X"0793F6F6";
				when "0001101101111"  => dbus <= X"00230300";
				when "0001101110000"  => dbus <= X"079300F5";
				when "0001101110001"  => dbus <= X"00A30780";
				when "0001101110010"  => dbus <= X"050900F5";
				when "0001101110011"  => dbus <= X"0785B795";
				when "0001101110100"  => dbus <= X"FFC78FA3";
				when "0001101110101"  => dbus <= X"40F60733";
				when "0001101110110"  => dbus <= X"FEE04BE3";
				when "0001101110111"  => dbus <= X"D36387B6";
				when "0001101111000"  => dbus <= X"47810006";
				when "0001101111001"  => dbus <= X"953E16FD";
				when "0001101111010"  => dbus <= X"B7A98E9D";
				when "0001101111011"  => dbus <= X"063387AA";
				when "0001101111100"  => dbus <= X"B7CD00D5";
				when "0001101111101"  => dbus <= X"0FA30505";
				when "0001101111110"  => dbus <= X"87B3FEE5";
				when "0001101111111"  => dbus <= X"4BE340A5";
				when "0001110000000"  => dbus <= X"87C2FEF8";
				when "0001110000001"  => dbus <= X"567D872A";
				when "0001110000010"  => dbus <= X"936317FD";
				when "0001110000011"  => dbus <= X"982A02C7";
				when "0001110000100"  => dbus <= X"05B38742";
				when "0001110000101"  => dbus <= X"051300D8";
				when "0001110000110"  => dbus <= X"86330200";
				when "0001110000111"  => dbus <= X"416340E5";
				when "0001110001000"  => dbus <= X"D36302C0";
				when "0001110001001"  => dbus <= X"46810006";
				when "0001110001010"  => dbus <= X"00D80533";
				when "0001110001011"  => dbus <= X"80826161";
				when "0001110001100"  => dbus <= X"95BE006C";
				when "0001110001101"  => dbus <= X"0005C583";
				when "0001110001110"  => dbus <= X"0FA30705";
				when "0001110001111"  => dbus <= X"B7E9FEB7";
				when "0001110010000"  => dbus <= X"0FA30705";
				when "0001110010001"  => dbus <= X"BFD1FEA7";
				when "0001110010010"  => dbus <= X"800007B7";
				when "0001110010011"  => dbus <= X"08A78023";
				when "0001110010100"  => dbus <= X"71498082";
				when "0001110010101"  => dbus <= X"14912223";
				when "0001110010110"  => dbus <= X"15212023";
				when "0001110010111"  => dbus <= X"13512A23";
				when "0001110011000"  => dbus <= X"14B12A23";
				when "0001110011001"  => dbus <= X"17012423";
				when "0001110011010"  => dbus <= X"08130ACC";
				when "0001110011011"  => dbus <= X"24B70201";
				when "0001110011100"  => dbus <= X"2AB74000";
				when "0001110011101"  => dbus <= X"29374000";
				when "0001110011110"  => dbus <= X"24234000";
				when "0001110011111"  => dbus <= X"2E231481";
				when "0001110100000"  => dbus <= X"26231331";
				when "0001110100001"  => dbus <= X"2C231411";
				when "0001110100010"  => dbus <= X"28231341";
				when "0001110100011"  => dbus <= X"26231361";
				when "0001110100100"  => dbus <= X"842A1371";
				when "0001110100101"  => dbus <= X"14C12C23";
				when "0001110100110"  => dbus <= X"14D12E23";
				when "0001110100111"  => dbus <= X"16E12023";
				when "0001110101000"  => dbus <= X"16F12223";
				when "0001110101001"  => dbus <= X"17112623";
				when "0001110101010"  => dbus <= X"89C2C22E";
				when "0001110101011"  => dbus <= X"15048493";
				when "0001110101100"  => dbus <= X"100A8A93";
				when "0001110101101"  => dbus <= X"12890913";
				when "0001110101110"  => dbus <= X"00044783";
				when "0001110101111"  => dbus <= X"0023E3A1";
				when "0001110110000"  => dbus <= X"45010008";
				when "0001110110001"  => dbus <= X"80000737";
				when "0001110110010"  => dbus <= X"00A987B3";
				when "0001110110011"  => dbus <= X"0007C783";
				when "0001110110100"  => dbus <= X"4A079763";
				when "0001110110101"  => dbus <= X"14C12083";
				when "0001110110110"  => dbus <= X"14812403";
				when "0001110110111"  => dbus <= X"14412483";
				when "0001110111000"  => dbus <= X"14012903";
				when "0001110111001"  => dbus <= X"13C12983";
				when "0001110111010"  => dbus <= X"13812A03";
				when "0001110111011"  => dbus <= X"13412A83";
				when "0001110111100"  => dbus <= X"13012B03";
				when "0001110111101"  => dbus <= X"12C12B83";
				when "0001110111110"  => dbus <= X"80826175";
				when "0001110111111"  => dbus <= X"02500713";
				when "0001111000000"  => dbus <= X"00E78863";
				when "0001111000001"  => dbus <= X"00180513";
				when "0001111000010"  => dbus <= X"00F80023";
				when "0001111000011"  => dbus <= X"A42D8A2E";
				when "0001111000100"  => dbus <= X"06934781";
				when "0001111000101"  => dbus <= X"051302B0";
				when "0001111000110"  => dbus <= X"089302D0";
				when "0001111000111"  => dbus <= X"03130300";
				when "0001111001000"  => dbus <= X"0E130200";
				when "0001111001001"  => dbus <= X"A8190230";
				when "0001111001010"  => dbus <= X"00A70763";
				when "0001111001011"  => dbus <= X"03171463";
				when "0001111001100"  => dbus <= X"0017E793";
				when "0001111001101"  => dbus <= X"E793A019";
				when "0001111001110"  => dbus <= X"84320107";
				when "0001111001111"  => dbus <= X"00144703";
				when "0001111010000"  => dbus <= X"00140613";
				when "0001111010001"  => dbus <= X"02D70363";
				when "0001111010010"  => dbus <= X"FEE6E0E3";
				when "0001111010011"  => dbus <= X"02670263";
				when "0001111010100"  => dbus <= X"03C70363";
				when "0001111010101"  => dbus <= X"FD070693";
				when "0001111010110"  => dbus <= X"0FF6F693";
				when "0001111010111"  => dbus <= X"62634525";
				when "0001111011000"  => dbus <= X"468106D5";
				when "0001111011001"  => dbus <= X"432948A5";
				when "0001111011010"  => dbus <= X"E793A005";
				when "0001111011011"  => dbus <= X"B7F10047";
				when "0001111011100"  => dbus <= X"0087E793";
				when "0001111011101"  => dbus <= X"E793B7D9";
				when "0001111011110"  => dbus <= X"B7C10207";
				when "0001111011111"  => dbus <= X"026686B3";
				when "0001111100000"  => dbus <= X"96AA0605";
				when "0001111100001"  => dbus <= X"FD068693";
				when "0001111100010"  => dbus <= X"00064503";
				when "0001111100011"  => dbus <= X"FD050713";
				when "0001111100100"  => dbus <= X"0FF77713";
				when "0001111100101"  => dbus <= X"FEE8F4E3";
				when "0001111100110"  => dbus <= X"00064503";
				when "0001111100111"  => dbus <= X"02E00713";
				when "0001111101000"  => dbus <= X"0CE51E63";
				when "0001111101001"  => dbus <= X"00164503";
				when "0001111101010"  => dbus <= X"041348A5";
				when "0001111101011"  => dbus <= X"07130016";
				when "0001111101100"  => dbus <= X"7713FD05";
				when "0001111101101"  => dbus <= X"E4630FF7";
				when "0001111101110"  => dbus <= X"47010AE8";
				when "0001111101111"  => dbus <= X"432948A5";
				when "0001111110000"  => dbus <= X"0513A03D";
				when "0001111110001"  => dbus <= X"56FD02A0";
				when "0001111110010"  => dbus <= X"FCA718E3";
				when "0001111110011"  => dbus <= X"06134194";
				when "0001111110100"  => dbus <= X"05910024";
				when "0001111110101"  => dbus <= X"FC06D2E3";
				when "0001111110110"  => dbus <= X"40D006B3";
				when "0001111110111"  => dbus <= X"0107E793";
				when "0001111111000"  => dbus <= X"0733BF65";
				when "0001111111001"  => dbus <= X"04050267";
				when "0001111111010"  => dbus <= X"0713972A";
				when "0001111111011"  => dbus <= X"4503FD07";
				when "0001111111100"  => dbus <= X"06130004";
				when "0001111111101"  => dbus <= X"7613FD05";
				when "0001111111110"  => dbus <= X"F4E30FF6";
				when "0001111111111"  => dbus <= X"4603FEC8";
				when "0010000000000"  => dbus <= X"05130004";
				when "0010000000001"  => dbus <= X"58FD04C0";
				when "0010000000010"  => dbus <= X"0DF67313";
				when "0010000000011"  => dbus <= X"00A31463";
				when "0010000000100"  => dbus <= X"040588B2";
				when "0010000000101"  => dbus <= X"00044503";
				when "0010000000110"  => dbus <= X"06900613";
				when "0010000000111"  => dbus <= X"06C50B63";
				when "0010000001000"  => dbus <= X"08A66163";
				when "0010000001001"  => dbus <= X"06100613";
				when "0010000001010"  => dbus <= X"18C50D63";
				when "0010000001011"  => dbus <= X"04A66B63";
				when "0010000001100"  => dbus <= X"04100613";
				when "0010000001101"  => dbus <= X"18C50563";
				when "0010000001110"  => dbus <= X"05800613";
				when "0010000001111"  => dbus <= X"32C50463";
				when "0010000010000"  => dbus <= X"02500793";
				when "0010000010001"  => dbus <= X"00F50563";
				when "0010000010010"  => dbus <= X"00F80023";
				when "0010000010011"  => dbus <= X"47830805";
				when "0010000010100"  => dbus <= X"99E30004";
				when "0010000010101"  => dbus <= X"147DEA07";
				when "0010000010110"  => dbus <= X"85428A2E";
				when "0010000010111"  => dbus <= X"0893A8F1";
				when "0010000011000"  => dbus <= X"470102A0";
				when "0010000011001"  => dbus <= X"F9151DE3";
				when "0010000011010"  => dbus <= X"04134198";
				when "0010000011011"  => dbus <= X"86130026";
				when "0010000011100"  => dbus <= X"53630045";
				when "0010000011101"  => dbus <= X"47010007";
				when "0010000011110"  => dbus <= X"B75185B2";
				when "0010000011111"  => dbus <= X"577D8432";
				when "0010000100000"  => dbus <= X"0613BFBD";
				when "0010000100001"  => dbus <= X"03630630";
				when "0010000100010"  => dbus <= X"061306C5";
				when "0010000100011"  => dbus <= X"19E30640";
				when "0010000100100"  => dbus <= X"0613FAC5";
				when "0010000100101"  => dbus <= X"E79306C0";
				when "0010000100110"  => dbus <= X"9B630027";
				when "0010000100111"  => dbus <= X"46292CC8";
				when "0010000101000"  => dbus <= X"0613A099";
				when "0010000101001"  => dbus <= X"01630730";
				when "0010000101010"  => dbus <= X"65630AC5";
				when "0010000101011"  => dbus <= X"061302A6";
				when "0010000101100"  => dbus <= X"0D6306F0";
				when "0010000101101"  => dbus <= X"06132AC5";
				when "0010000101110"  => dbus <= X"13E30700";
				when "0010000101111"  => dbus <= X"567DF8C5";
				when "0010000110000"  => dbus <= X"00C69563";
				when "0010000110001"  => dbus <= X"0017E793";
				when "0010000110010"  => dbus <= X"8A1346A1";
				when "0010000110011"  => dbus <= X"46410045";
				when "0010000110100"  => dbus <= X"A45D418C";
				when "0010000110101"  => dbus <= X"07500613";
				when "0010000110110"  => dbus <= X"FCC503E3";
				when "0010000110111"  => dbus <= X"07800313";
				when "0010000111000"  => dbus <= X"1FE34641";
				when "0010000111001"  => dbus <= X"8A13F465";
				when "0010000111010"  => dbus <= X"B7DD0045";
				when "0010000111011"  => dbus <= X"E79D8BC1";
				when "0010000111100"  => dbus <= X"00D80633";
				when "0010000111101"  => dbus <= X"02000513";
				when "0010000111110"  => dbus <= X"8FA3A021";
				when "0010000111111"  => dbus <= X"883EFEA7";
				when "0010001000000"  => dbus <= X"00180793";
				when "0010001000001"  => dbus <= X"40F60733";
				when "0010001000010"  => dbus <= X"FEE049E3";
				when "0010001000011"  => dbus <= X"FFF68793";
				when "0010001000100"  => dbus <= X"00D04363";
				when "0010001000101"  => dbus <= X"86B34685";
				when "0010001000110"  => dbus <= X"068540D7";
				when "0010001000111"  => dbus <= X"8A13419C";
				when "0010001001000"  => dbus <= X"05130045";
				when "0010001001001"  => dbus <= X"00230018";
				when "0010001001010"  => dbus <= X"96C200F8";
				when "0010001001011"  => dbus <= X"02000713";
				when "0010001001100"  => dbus <= X"40A687B3";
				when "0010001001101"  => dbus <= X"00F04663";
				when "0010001001110"  => dbus <= X"85D20405";
				when "0010001001111"  => dbus <= X"BBAD882A";
				when "0010001010000"  => dbus <= X"0FA30505";
				when "0010001010001"  => dbus <= X"B7EDFEE5";
				when "0010001010010"  => dbus <= X"00458A13";
				when "0010001010011"  => dbus <= X"E191418C";
				when "0010001010100"  => dbus <= X"972E85A6";
				when "0010001010101"  => dbus <= X"4503862E";
				when "0010001010110"  => dbus <= X"C1190006";
				when "0010001010111"  => dbus <= X"02E61B63";
				when "0010001011000"  => dbus <= X"07338BC1";
				when "0010001011001"  => dbus <= X"061340B6";
				when "0010001011010"  => dbus <= X"CB950200";
				when "0010001011011"  => dbus <= X"CE634781";
				when "0010001011100"  => dbus <= X"853A02E7";
				when "0010001011101"  => dbus <= X"00075363";
				when "0010001011110"  => dbus <= X"95424501";
				when "0010001011111"  => dbus <= X"061396AA";
				when "0010001100000"  => dbus <= X"87B30200";
				when "0010001100001"  => dbus <= X"59E340A6";
				when "0010001100010"  => dbus <= X"0505FAF7";
				when "0010001100011"  => dbus <= X"FEC50FA3";
				when "0010001100100"  => dbus <= X"0605BFCD";
				when "0010001100101"  => dbus <= X"0805B7C9";
				when "0010001100110"  => dbus <= X"FEC80FA3";
				when "0010001100111"  => dbus <= X"879386BE";
				when "0010001101000"  => dbus <= X"4AE3FFF6";
				when "0010001101001"  => dbus <= X"86BEFED7";
				when "0010001101010"  => dbus <= X"8633B7D1";
				when "0010001101011"  => dbus <= X"450300F5";
				when "0010001101100"  => dbus <= X"06330006";
				when "0010001101101"  => dbus <= X"078500F8";
				when "0010001101110"  => dbus <= X"00A60023";
				when "0010001101111"  => dbus <= X"E793BF4D";
				when "0010001110000"  => dbus <= X"07130407";
				when "0010001110001"  => dbus <= X"AE0306C0";
				when "0010001110010"  => dbus <= X"8A130005";
				when "0010001110011"  => dbus <= X"91630045";
				when "0010001110100"  => dbus <= X"F71310E8";
				when "0010001110101"  => dbus <= X"85560407";
				when "0010001110110"  => dbus <= X"854AC311";
				when "0010001110111"  => dbus <= X"45810038";
				when "0010001111000"  => dbus <= X"4E99833A";
				when "0010001111001"  => dbus <= X"03A00F13";
				when "0010001111010"  => dbus <= X"00BE0633";
				when "0010001111011"  => dbus <= X"00064603";
				when "0010001111100"  => dbus <= X"070D0585";
				when "0010001111101"  => dbus <= X"00465893";
				when "0010001111110"  => dbus <= X"98AA8A3D";
				when "0010001111111"  => dbus <= X"C883962A";
				when "0010010000000"  => dbus <= X"46030008";
				when "0010010000001"  => dbus <= X"0EA30006";
				when "0010010000010"  => dbus <= X"0F23FF17";
				when "0010010000011"  => dbus <= X"9763FEC7";
				when "0010010000100"  => dbus <= X"8BC105D5";
				when "0010010000101"  => dbus <= X"4645EB99";
				when "0010010000110"  => dbus <= X"02000593";
				when "0010010000111"  => dbus <= X"FFF68793";
				when "0010010001000"  => dbus <= X"00180713";
				when "0010010001001"  => dbus <= X"02D64F63";
				when "0010010001010"  => dbus <= X"478186BE";
				when "0010010001011"  => dbus <= X"05B34745";
				when "0010010001100"  => dbus <= X"C58300F3";
				when "0010010001101"  => dbus <= X"06330005";
				when "0010010001110"  => dbus <= X"078500F8";
				when "0010010001111"  => dbus <= X"00B60023";
				when "0010010010000"  => dbus <= X"FEE797E3";
				when "0010010010001"  => dbus <= X"01180513";
				when "0010010010010"  => dbus <= X"071347C5";
				when "0010010010011"  => dbus <= X"D5E30200";
				when "0010010010100"  => dbus <= X"0505EED7";
				when "0010010010101"  => dbus <= X"FEE50FA3";
				when "0010010010110"  => dbus <= X"BFD516FD";
				when "0010010010111"  => dbus <= X"FFE70FA3";
				when "0010010011000"  => dbus <= X"0FA3B761";
				when "0010010011001"  => dbus <= X"86BEFEB7";
				when "0010010011010"  => dbus <= X"BF4D883A";
				when "0010010011011"  => dbus <= X"05931218";
				when "0010010011100"  => dbus <= X"963A0016";
				when "0010010011101"  => dbus <= X"EF660423";
				when "0010010011110"  => dbus <= X"00AE0733";
				when "0010010011111"  => dbus <= X"00074703";
				when "0010010100000"  => dbus <= X"12010313";
				when "0010010100001"  => dbus <= X"00158613";
				when "0010010100010"  => dbus <= X"E32D932E";
				when "0010010100011"  => dbus <= X"EE730423";
				when "0010010100100"  => dbus <= X"1DE30505";
				when "0010010100101"  => dbus <= X"8BC1FDE5";
				when "0010010100110"  => dbus <= X"02000593";
				when "0010010100111"  => dbus <= X"4781CFC5";
				when "0010010101000"  => dbus <= X"95BE002C";
				when "0010010101001"  => dbus <= X"0005C583";
				when "0010010101010"  => dbus <= X"00F80733";
				when "0010010101011"  => dbus <= X"00230785";
				when "0010010101100"  => dbus <= X"97E300B7";
				when "0010010101101"  => dbus <= X"0533FEC7";
				when "0010010101110"  => dbus <= X"96AA00C8";
				when "0010010101111"  => dbus <= X"02000713";
				when "0010010110000"  => dbus <= X"40A687B3";
				when "0010010110001"  => dbus <= X"E6F65AE3";
				when "0010010110010"  => dbus <= X"0FA30505";
				when "0010010110011"  => dbus <= X"BFCDFEE5";
				when "0010010110100"  => dbus <= X"45814501";
				when "0010010110101"  => dbus <= X"06300F93";
				when "0010010110110"  => dbus <= X"48A942A5";
				when "0010010110111"  => dbus <= X"06400E93";
				when "0010010111000"  => dbus <= X"03000393";
				when "0010010111001"  => dbus <= X"0B134F11";
				when "0010010111010"  => dbus <= X"B77902E0";
				when "0010010111011"  => dbus <= X"04EFD363";
				when "0010010111100"  => dbus <= X"03D74BB3";
				when "0010010111101"  => dbus <= X"67330589";
				when "0010010111110"  => dbus <= X"9BD603D7";
				when "0010010111111"  => dbus <= X"000BCB83";
				when "0010011000000"  => dbus <= X"EF730423";
				when "0010011000001"  => dbus <= X"12010313";
				when "0010011000010"  => dbus <= X"4333961A";
				when "0010011000011"  => dbus <= X"67330317";
				when "0010011000100"  => dbus <= X"93560317";
				when "0010011000101"  => dbus <= X"00034303";
				when "0010011000110"  => dbus <= X"EE660423";
				when "0010011000111"  => dbus <= X"47039756";
				when "0010011001000"  => dbus <= X"03130007";
				when "0010011001001"  => dbus <= X"86131201";
				when "0010011001010"  => dbus <= X"959A0015";
				when "0010011001011"  => dbus <= X"EEE58423";
				when "0010011001100"  => dbus <= X"D5E3B785";
				when "0010011001101"  => dbus <= X"45B3FEE2";
				when "0010011001110"  => dbus <= X"95D60317";
				when "0010011001111"  => dbus <= X"0005C583";
				when "0010011010000"  => dbus <= X"03176733";
				when "0010011010001"  => dbus <= X"EEB30423";
				when "0010011010010"  => dbus <= X"BFC985B2";
				when "0010011010011"  => dbus <= X"FEB70FA3";
				when "0010011010100"  => dbus <= X"883A86BE";
				when "0010011010101"  => dbus <= X"FFF68793";
				when "0010011010110"  => dbus <= X"00180713";
				when "0010011010111"  => dbus <= X"FED648E3";
				when "0010011011000"  => dbus <= X"BF3586BE";
				when "0010011011001"  => dbus <= X"0407E793";
				when "0010011011010"  => dbus <= X"BBB54641";
				when "0010011011011"  => dbus <= X"BBA54621";
				when "0010011011100"  => dbus <= X"00458A13";
				when "0010011011101"  => dbus <= X"4629418C";
				when "0010011011110"  => dbus <= X"3A398542";
				when "0010011011111"  => dbus <= X"0023BB75";
				when "0010011100000"  => dbus <= X"050508F7";
				when "0010011100001"  => dbus <= X"27F3B691";
				when "0010011100010"  => dbus <= X"2573C810";
				when "0010011100011"  => dbus <= X"25F3C010";
				when "0010011100100"  => dbus <= X"9AE3C810";
				when "0010011100101"  => dbus <= X"8082FEF5";
				when "0010011100110"  => dbus <= X"C4221141";
				when "0010011100111"  => dbus <= X"C606C226";
				when "0010011101000"  => dbus <= X"84AE842A";
				when "0010011101001"  => dbus <= X"07B337CD";
				when "0010011101010"  => dbus <= X"B5330085";
				when "0010011101011"  => dbus <= X"95A600A7";
				when "0010011101100"  => dbus <= X"577D952E";
				when "0010011101101"  => dbus <= X"88371073";
				when "0010011101110"  => dbus <= X"80379073";
				when "0010011101111"  => dbus <= X"88351073";
				when "0010011110000"  => dbus <= X"442240B2";
				when "0010011110001"  => dbus <= X"01414492";
				when "0010011110010"  => dbus <= X"47818082";
				when "0010011110011"  => dbus <= X"00C79363";
				when "0010011110100"  => dbus <= X"87338082";
				when "0010011110101"  => dbus <= X"468300F5";
				when "0010011110110"  => dbus <= X"07330007";
				when "0010011110111"  => dbus <= X"078500F5";
				when "0010011111000"  => dbus <= X"00D70023";
				when "0010011111001"  => dbus <= X"07B7B7E5";
				when "0010011111010"  => dbus <= X"80238000";
				when "0010011111011"  => dbus <= X"808208A7";
				when "0010011111100"  => dbus <= X"80000737";
				when "0010011111101"  => dbus <= X"00054783";
				when "0010011111110"  => dbus <= X"8082E391";
				when "0010011111111"  => dbus <= X"00230505";
				when "0010100000000"  => dbus <= X"BFCD08F7";
				when "0010100000001"  => dbus <= X"005C1141";
				when "0010100000010"  => dbus <= X"472986BE";
				when "0010100000011"  => dbus <= X"8163E115";
				when "0010100000100"  => dbus <= X"063702D7";
				when "0010100000101"  => dbus <= X"17FD8000";
				when "0010100000110"  => dbus <= X"0007C703";
				when "0010100000111"  => dbus <= X"03070713";
				when "0010100001000"  => dbus <= X"0FF77713";
				when "0010100001001"  => dbus <= X"08E60023";
				when "0010100001010"  => dbus <= X"FED797E3";
				when "0010100001011"  => dbus <= X"80820141";
				when "0010100001100"  => dbus <= X"02E57633";
				when "0010100001101"  => dbus <= X"8FA30785";
				when "0010100001110"  => dbus <= X"5533FEC7";
				when "0010100001111"  => dbus <= X"B7F902E5";
				when "0010100010000"  => dbus <= X"273715FD";
				when "0010100010001"  => dbus <= X"058A4000";
				when "0010100010010"  => dbus <= X"15870713";
				when "0010100010011"  => dbus <= X"800006B7";
				when "0010100010100"  => dbus <= X"0005D363";
				when "0010100010101"  => dbus <= X"57B38082";
				when "0010100010110"  => dbus <= X"8BBD00B5";
				when "0010100010111"  => dbus <= X"C78397BA";
				when "0010100011000"  => dbus <= X"15F10007";
				when "0010100011001"  => dbus <= X"08F68023";
				when "0010100011010"  => dbus <= X"0737B7E5";
				when "0010100011011"  => dbus <= X"475C8000";
				when "0010100011100"  => dbus <= X"DFF58B85";
				when "0010100011101"  => dbus <= X"8082C348";
				when "0010100011110"  => dbus <= X"80000737";
				when "0010100011111"  => dbus <= X"8B89475C";
				when "0010100100000"  => dbus <= X"4308DFF5";
				when "0010100100001"  => dbus <= X"0FF57513";
				when "0010100100010"  => dbus <= X"07378082";
				when "0010100100011"  => dbus <= X"4F5C8000";
				when "0010100100100"  => dbus <= X"DFF58B85";
				when "0010100100101"  => dbus <= X"8082CB48";
				when "0010100100110"  => dbus <= X"80000737";
				when "0010100100111"  => dbus <= X"8B894F5C";
				when "0010100101000"  => dbus <= X"4B08DFF5";
				when "0010100101001"  => dbus <= X"0FF57513";
				when "0010100101010"  => dbus <= X"11418082";
				when "0010100101011"  => dbus <= X"C606C422";
				when "0010100101100"  => dbus <= X"4503842A";
				when "0010100101101"  => dbus <= X"E5090004";
				when "0010100101110"  => dbus <= X"442240B2";
				when "0010100101111"  => dbus <= X"80820141";
				when "0010100110000"  => dbus <= X"37650405";
				when "0010100110001"  => dbus <= X"1141B7FD";
				when "0010100110010"  => dbus <= X"C606C422";
				when "0010100110011"  => dbus <= X"4503842A";
				when "0010100110100"  => dbus <= X"E5090004";
				when "0010100110101"  => dbus <= X"442240B2";
				when "0010100110110"  => dbus <= X"80820141";
				when "0010100110111"  => dbus <= X"37750405";
				when "0010100111000"  => dbus <= X"7159B7FD";
				when "0010100111001"  => dbus <= X"6705D686";
				when "0010100111010"  => dbus <= X"D2A6D4A2";
				when "0010100111011"  => dbus <= X"CECED0CA";
				when "0010100111100"  => dbus <= X"CAD6CCD2";
				when "0010100111101"  => dbus <= X"C6DEC8DA";
				when "0010100111110"  => dbus <= X"C2E6C4E2";
				when "0010100111111"  => dbus <= X"81010113";
				when "0010101000000"  => dbus <= X"07930814";
				when "0010101000001"  => dbus <= X"75FD8207";
				when "0010101000010"  => dbus <= X"861397B6";
				when "0010101000011"  => dbus <= X"963E7E85";
				when "0010101000100"  => dbus <= X"82070793";
				when "0010101000101"  => dbus <= X"859397B6";
				when "0010101000110"  => dbus <= X"95BE7E45";
				when "0010101000111"  => dbus <= X"05E10513";
				when "0010101001000"  => dbus <= X"F0EFCA02";
				when "0010101001001"  => dbus <= X"4505BCEF";
				when "0010101001010"  => dbus <= X"ECAFF0EF";
				when "0010101001011"  => dbus <= X"00A11E23";
				when "0010101001100"  => dbus <= X"F0EF4509";
				when "0010101001101"  => dbus <= X"1F23EC0F";
				when "0010101001110"  => dbus <= X"450D00A1";
				when "0010101001111"  => dbus <= X"EB6FF0EF";
				when "0010101010000"  => dbus <= X"02A11023";
				when "0010101010001"  => dbus <= X"F0EF4511";
				when "0010101010010"  => dbus <= X"DC2AEACF";
				when "0010101010011"  => dbus <= X"F0EF4515";
				when "0010101010100"  => dbus <= X"0063EA4F";
				when "0010101010101"  => dbus <= X"DE2A3805";
				when "0010101010110"  => dbus <= X"07136705";
				when "0010101010111"  => dbus <= X"08148207";
				when "0010101011000"  => dbus <= X"973677FD";
				when "0010101011001"  => dbus <= X"C63E97BA";
				when "0010101011010"  => dbus <= X"7EC7A783";
				when "0010101011011"  => dbus <= X"47B2EB91";
				when "0010101011100"  => dbus <= X"7F079783";
				when "0010101011101"  => dbus <= X"4732E3B1";
				when "0010101011110"  => dbus <= X"06600793";
				when "0010101011111"  => dbus <= X"7EF71823";
				when "0010101100000"  => dbus <= X"07136705";
				when "0010101100001"  => dbus <= X"08148207";
				when "0010101100010"  => dbus <= X"77FD9736";
				when "0010101100011"  => dbus <= X"A70397BA";
				when "0010101100100"  => dbus <= X"C63E7EC7";
				when "0010101100101"  => dbus <= X"11634785";
				when "0010101100110"  => dbus <= X"47B202F7";
				when "0010101100111"  => dbus <= X"7F079783";
				when "0010101101000"  => dbus <= X"4732EF81";
				when "0010101101001"  => dbus <= X"341537B7";
				when "0010101101010"  => dbus <= X"41578793";
				when "0010101101011"  => dbus <= X"7EF72623";
				when "0010101101100"  => dbus <= X"06600793";
				when "0010101101101"  => dbus <= X"7EF71823";
				when "0010101101110"  => dbus <= X"08146705";
				when "0010101101111"  => dbus <= X"82070713";
				when "0010101110000"  => dbus <= X"77FD9736";
				when "0010101110001"  => dbus <= X"C63E97BA";
				when "0010101110010"  => dbus <= X"473256F2";
				when "0010101110011"  => dbus <= X"F313109C";
				when "0010101110100"  => dbus <= X"2A230016";
				when "0010101110101"  => dbus <= X"1E237EF7";
				when "0010101110110"  => dbus <= X"F7930401";
				when "0010101110111"  => dbus <= X"851A0026";
				when "0010101111000"  => dbus <= X"0513C399";
				when "0010101111001"  => dbus <= X"F7930013";
				when "0010101111010"  => dbus <= X"C7810046";
				when "0010101111011"  => dbus <= X"05420505";
				when "0010101111100"  => dbus <= X"07938141";
				when "0010101111101"  => dbus <= X"D5337D00";
				when "0010101111110"  => dbus <= X"648502A7";
				when "0010101111111"  => dbus <= X"0813767D";
				when "0010110000000"  => dbus <= X"84130101";
				when "0010110000001"  => dbus <= X"05938204";
				when "0010110000010"  => dbus <= X"94427EC6";
				when "0010110000011"  => dbus <= X"841395A2";
				when "0010110000100"  => dbus <= X"94428204";
				when "0010110000101"  => dbus <= X"47014781";
				when "0010110000110"  => dbus <= X"96224E85";
				when "0010110000111"  => dbus <= X"DA2A4E0D";
				when "0010110001000"  => dbus <= X"00FE9833";
				when "0010110001001"  => dbus <= X"00D87833";
				when "0010110001010"  => dbus <= X"00080F63";
				when "0010110001011"  => dbus <= X"02A70F33";
				when "0010110001100"  => dbus <= X"7F462883";
				when "0010110001101"  => dbus <= X"00279813";
				when "0010110001110"  => dbus <= X"982E0705";
				when "0010110001111"  => dbus <= X"83410742";
				when "0010110010000"  => dbus <= X"262398FA";
				when "0010110010001"  => dbus <= X"07850118";
				when "0010110010010"  => dbus <= X"FDC79CE3";
				when "0010110010011"  => dbus <= X"02030163";
				when "0010110010100"  => dbus <= X"08146705";
				when "0010110010101"  => dbus <= X"82070713";
				when "0010110010110"  => dbus <= X"77FD9736";
				when "0010110010111"  => dbus <= X"960397BA";
				when "0010110011000"  => dbus <= X"A5837EC7";
				when "0010110011001"  => dbus <= X"C63E7F87";
				when "0010110011010"  => dbus <= X"E37FE0EF";
				when "0010110011011"  => dbus <= X"6705C0AA";
				when "0010110011100"  => dbus <= X"82070713";
				when "0010110011101"  => dbus <= X"77FD0814";
				when "0010110011110"  => dbus <= X"97BA9736";
				when "0010110011111"  => dbus <= X"57F2C63E";
				when "0010110100000"  => dbus <= X"CF998B89";
				when "0010110100001"  => dbus <= X"473247B2";
				when "0010110100010"  => dbus <= X"97835552";
				when "0010110100011"  => dbus <= X"16037EE7";
				when "0010110100100"  => dbus <= X"25837EC7";
				when "0010110100101"  => dbus <= X"07C27FC7";
				when "0010110100110"  => dbus <= X"8E5D00D4";
				when "0010110100111"  => dbus <= X"EFBFE0EF";
				when "0010110101000"  => dbus <= X"777D57F2";
				when "0010110101001"  => dbus <= X"CF918B91";
				when "0010110101010"  => dbus <= X"87936785";
				when "0010110101011"  => dbus <= X"08148207";
				when "0010110101100"  => dbus <= X"97BA97B6";
				when "0010110101101"  => dbus <= X"95835642";
				when "0010110101110"  => dbus <= X"55527EC7";
				when "0010110101111"  => dbus <= X"F0EFC63E";
				when "0010110110000"  => dbus <= X"57E2A58F";
				when "0010110110001"  => dbus <= X"4785E7A1";
				when "0010110110010"  => dbus <= X"6785DC3E";
				when "0010110110011"  => dbus <= X"879374FD";
				when "0010110110100"  => dbus <= X"08188207";
				when "0010110110101"  => dbus <= X"7EC48493";
				when "0010110110110"  => dbus <= X"442997BA";
				when "0010110110111"  => dbus <= X"57E294BE";
				when "0010110111000"  => dbus <= X"028787B3";
				when "0010110111001"  => dbus <= X"F0EFDC3E";
				when "0010110111010"  => dbus <= X"85269C0F";
				when "0010110111011"  => dbus <= X"975FE0EF";
				when "0010110111100"  => dbus <= X"9D0FF0EF";
				when "0010110111101"  => dbus <= X"9E6FF0EF";
				when "0010110111110"  => dbus <= X"9EEFF0EF";
				when "0010110111111"  => dbus <= X"5433D16D";
				when "0010111000000"  => dbus <= X"556202A4";
				when "0010111000001"  => dbus <= X"04330405";
				when "0010111000010"  => dbus <= X"DC2202A4";
				when "0010111000011"  => dbus <= X"99AFF0EF";
				when "0010111000100"  => dbus <= X"08186485";
				when "0010111000101"  => dbus <= X"8793747D";
				when "0010111000110"  => dbus <= X"97BA8204";
				when "0010111000111"  => dbus <= X"7EC40513";
				when "0010111001000"  => dbus <= X"E0EF953E";
				when "0010111001001"  => dbus <= X"F0EF93FF";
				when "0010111001010"  => dbus <= X"F0EF99AF";
				when "0010111001011"  => dbus <= X"08189B0F";
				when "0010111001100"  => dbus <= X"82048793";
				when "0010111001101"  => dbus <= X"97A297BA";
				when "0010111001110"  => dbus <= X"95038B2A";
				when "0010111001111"  => dbus <= X"45817EC7";
				when "0010111010000"  => dbus <= X"F0EFC63E";
				when "0010111010001"  => dbus <= X"47B2D4CF";
				when "0010111010010"  => dbus <= X"950385AA";
				when "0010111010011"  => dbus <= X"F0EF7EE7";
				when "0010111010100"  => dbus <= X"47B2D40F";
				when "0010111010101"  => dbus <= X"950385AA";
				when "0010111010110"  => dbus <= X"F0EF7F07";
				when "0010111010111"  => dbus <= X"85AAD34F";
				when "0010111011000"  => dbus <= X"03411503";
				when "0010111011001"  => dbus <= X"D2AFF0EF";
				when "0010111011010"  => dbus <= X"879367A1";
				when "0010111011011"  => dbus <= X"89AAB057";
				when "0010111011100"  => dbus <= X"1CF50163";
				when "0010111011101"  => dbus <= X"16A7E263";
				when "0010111011110"  => dbus <= X"87936789";
				when "0010111011111"  => dbus <= X"0A638F27";
				when "0010111100000"  => dbus <= X"67951CF5";
				when "0010111100001"  => dbus <= X"EAF78793";
				when "0010111100010"  => dbus <= X"1AF50D63";
				when "0010111100011"  => dbus <= X"F0EF547D";
				when "0010111100100"  => dbus <= X"55D2D06F";
				when "0010111100101"  => dbus <= X"2537942A";
				when "0010111100110"  => dbus <= X"05134000";
				when "0010111100111"  => dbus <= X"F0EFD745";
				when "0010111101000"  => dbus <= X"2537EB4F";
				when "0010111101001"  => dbus <= X"85DA4000";
				when "0010111101010"  => dbus <= X"D8C50513";
				when "0010111101011"  => dbus <= X"EA6FF0EF";
				when "0010111101100"  => dbus <= X"F0EF855A";
				when "0010111101101"  => dbus <= X"85AA934F";
				when "0010111101110"  => dbus <= X"40002537";
				when "0010111101111"  => dbus <= X"DA450513";
				when "0010111110000"  => dbus <= X"E92FF0EF";
				when "0010111110001"  => dbus <= X"855A0442";
				when "0010111110010"  => dbus <= X"F0EF8041";
				when "0010111110011"  => dbus <= X"C10D91CF";
				when "0010111110100"  => dbus <= X"00C02583";
				when "0010111110101"  => dbus <= X"855A54E2";
				when "0010111110110"  => dbus <= X"02B484B3";
				when "0010111110111"  => dbus <= X"90AFF0EF";
				when "0010111111000"  => dbus <= X"02A4D5B3";
				when "0010111111001"  => dbus <= X"40002537";
				when "0010111111010"  => dbus <= X"DBC50513";
				when "0010111111011"  => dbus <= X"E66FF0EF";
				when "0010111111100"  => dbus <= X"F0EF855A";
				when "0010111111101"  => dbus <= X"47A58F4F";
				when "0010111111110"  => dbus <= X"24A7F163";
				when "0010111111111"  => dbus <= X"00C02783";
				when "0011000000000"  => dbus <= X"253755E2";
				when "0011000000001"  => dbus <= X"05134000";
				when "0011000000010"  => dbus <= X"85B3E145";
				when "0011000000011"  => dbus <= X"044202F5";
				when "0011000000100"  => dbus <= X"F0EF8441";
				when "0011000000101"  => dbus <= X"25B7E40F";
				when "0011000000110"  => dbus <= X"25374000";
				when "0011000000111"  => dbus <= X"85934000";
				when "0011000001000"  => dbus <= X"0513E2C5";
				when "0011000001001"  => dbus <= X"F0EFE385";
				when "0011000001010"  => dbus <= X"25B7E2CF";
				when "0011000001011"  => dbus <= X"25374000";
				when "0011000001100"  => dbus <= X"85934000";
				when "0011000001101"  => dbus <= X"0513E505";
				when "0011000001110"  => dbus <= X"F0EFE745";
				when "0011000001111"  => dbus <= X"25B7E18F";
				when "0011000010000"  => dbus <= X"25374000";
				when "0011000010001"  => dbus <= X"85934000";
				when "0011000010010"  => dbus <= X"0513E8C5";
				when "0011000010011"  => dbus <= X"F0EFE945";
				when "0011000010100"  => dbus <= X"2537E04F";
				when "0011000010101"  => dbus <= X"85CE4000";
				when "0011000010110"  => dbus <= X"EAC50513";
				when "0011000010111"  => dbus <= X"DF6FF0EF";
				when "0011000011000"  => dbus <= X"8B8557F2";
				when "0011000011001"  => dbus <= X"20079663";
				when "0011000011010"  => dbus <= X"8B8957F2";
				when "0011000011011"  => dbus <= X"24079363";
				when "0011000011100"  => dbus <= X"8B9157F2";
				when "0011000011101"  => dbus <= X"28079063";
				when "0011000011110"  => dbus <= X"87936785";
				when "0011000011111"  => dbus <= X"08188207";
				when "0011000100000"  => dbus <= X"97BA79FD";
				when "0011000100001"  => dbus <= X"99BE4481";
				when "0011000100010"  => dbus <= X"04400A13";
				when "0011000100011"  => dbus <= X"2B376A85";
				when "0011000100100"  => dbus <= X"27834000";
				when "0011000100101"  => dbus <= X"ED6300C0";
				when "0011000100110"  => dbus <= X"1A6326F4";
				when "0011000100111"  => dbus <= X"25372804";
				when "0011000101000"  => dbus <= X"05134000";
				when "0011000101001"  => dbus <= X"F0EFF385";
				when "0011000101010"  => dbus <= X"0513DACF";
				when "0011000101011"  => dbus <= X"F0EF05E1";
				when "0011000101100"  => dbus <= X"0113862F";
				when "0011000101101"  => dbus <= X"50B67F01";
				when "0011000101110"  => dbus <= X"54264501";
				when "0011000101111"  => dbus <= X"59065496";
				when "0011000110000"  => dbus <= X"4A6649F6";
				when "0011000110001"  => dbus <= X"4B464AD6";
				when "0011000110010"  => dbus <= X"4C264BB6";
				when "0011000110011"  => dbus <= X"61654C96";
				when "0011000110100"  => dbus <= X"479D8082";
				when "0011000110101"  => dbus <= X"B149DE3E";
				when "0011000110110"  => dbus <= X"879367A5";
				when "0011000110111"  => dbus <= X"0F63A027";
				when "0011000111000"  => dbus <= X"67BD00F5";
				when "0011000111001"  => dbus <= X"9F578793";
				when "0011000111010"  => dbus <= X"EAF512E3";
				when "0011000111011"  => dbus <= X"40002537";
				when "0011000111100"  => dbus <= X"C8450513";
				when "0011000111101"  => dbus <= X"D5EFF0EF";
				when "0011000111110"  => dbus <= X"A801478D";
				when "0011000111111"  => dbus <= X"40002537";
				when "0011001000000"  => dbus <= X"BF450513";
				when "0011001000001"  => dbus <= X"D4EFF0EF";
				when "0011001000010"  => dbus <= X"67054781";
				when "0011001000011"  => dbus <= X"82070713";
				when "0011001000100"  => dbus <= X"2A370814";
				when "0011001000101"  => dbus <= X"7BFD4000";
				when "0011001000110"  => dbus <= X"07869736";
				when "0011001000111"  => dbus <= X"B48A0A13";
				when "0011001001000"  => dbus <= X"44814401";
				when "0011001001001"  => dbus <= X"9A3E9BBA";
				when "0011001001010"  => dbus <= X"40002C37";
				when "0011001001011"  => dbus <= X"40002CB7";
				when "0011001001100"  => dbus <= X"2537A201";
				when "0011001001101"  => dbus <= X"05134000";
				when "0011001001110"  => dbus <= X"F0EFC245";
				when "0011001001111"  => dbus <= X"4785D18F";
				when "0011001010000"  => dbus <= X"2537B7E9";
				when "0011001010001"  => dbus <= X"05134000";
				when "0011001010010"  => dbus <= X"F0EFC505";
				when "0011001010011"  => dbus <= X"4789D08F";
				when "0011001010100"  => dbus <= X"2537BF6D";
				when "0011001010101"  => dbus <= X"05134000";
				when "0011001010110"  => dbus <= X"F0EFCB45";
				when "0011001010111"  => dbus <= X"4791CF8F";
				when "0011001011000"  => dbus <= X"0A93B76D";
				when "0011001011001"  => dbus <= X"8AB30440";
				when "0011001011010"  => dbus <= X"87B30354";
				when "0011001011011"  => dbus <= X"6A85015B";
				when "0011001011100"  => dbus <= X"A7839ABE";
				when "0011001011101"  => dbus <= X"962380CA";
				when "0011001011110"  => dbus <= X"8B85820A";
				when "0011001011111"  => dbus <= X"D603C38D";
				when "0011001100000"  => dbus <= X"5683826A";
				when "0011001100001"  => dbus <= X"0C63000A";
				when "0011001100010"  => dbus <= X"85A600D6";
				when "0011001100011"  => dbus <= X"CE0C0513";
				when "0011001100100"  => dbus <= X"CC2FF0EF";
				when "0011001100101"  => dbus <= X"82CAD783";
				when "0011001100110"  => dbus <= X"96230785";
				when "0011001100111"  => dbus <= X"0A9382FA";
				when "0011001101000"  => dbus <= X"8AB30440";
				when "0011001101001"  => dbus <= X"87B30354";
				when "0011001101010"  => dbus <= X"6A85015B";
				when "0011001101011"  => dbus <= X"A7839ABE";
				when "0011001101100"  => dbus <= X"8B8980CA";
				when "0011001101101"  => dbus <= X"D603C38D";
				when "0011001101110"  => dbus <= X"5683828A";
				when "0011001101111"  => dbus <= X"0C6300CA";
				when "0011001110000"  => dbus <= X"85A600D6";
				when "0011001110001"  => dbus <= X"D10C8513";
				when "0011001110010"  => dbus <= X"C8AFF0EF";
				when "0011001110011"  => dbus <= X"82CAD783";
				when "0011001110100"  => dbus <= X"96230785";
				when "0011001110101"  => dbus <= X"0A9382FA";
				when "0011001110110"  => dbus <= X"8AB30440";
				when "0011001110111"  => dbus <= X"87B30354";
				when "0011001111000"  => dbus <= X"6A85015B";
				when "0011001111001"  => dbus <= X"A7839ABE";
				when "0011001111010"  => dbus <= X"8B9180CA";
				when "0011001111011"  => dbus <= X"D603C39D";
				when "0011001111100"  => dbus <= X"568382AA";
				when "0011001111101"  => dbus <= X"0E63018A";
				when "0011001111110"  => dbus <= X"253700D6";
				when "0011001111111"  => dbus <= X"85A64000";
				when "0011010000000"  => dbus <= X"D4450513";
				when "0011010000001"  => dbus <= X"C4EFF0EF";
				when "0011010000010"  => dbus <= X"82CAD783";
				when "0011010000011"  => dbus <= X"96230785";
				when "0011010000100"  => dbus <= X"079382FA";
				when "0011010000101"  => dbus <= X"87B30440";
				when "0011010000110"  => dbus <= X"670502F4";
				when "0011010000111"  => dbus <= X"04C20485";
				when "0011010001000"  => dbus <= X"97DE80C1";
				when "0011010001001"  => dbus <= X"D50397BA";
				when "0011010001010"  => dbus <= X"942A82C7";
				when "0011010001011"  => dbus <= X"84410442";
				when "0011010001100"  => dbus <= X"00C02783";
				when "0011010001101"  => dbus <= X"F2F4E7E3";
				when "0011010001110"  => dbus <= X"2537BB99";
				when "0011010001111"  => dbus <= X"05134000";
				when "0011010010000"  => dbus <= X"F0EFDD45";
				when "0011010010001"  => dbus <= X"0405C10F";
				when "0011010010010"  => dbus <= X"87B3BB55";
				when "0011010010011"  => dbus <= X"85A60344";
				when "0011010010100"  => dbus <= X"05130485";
				when "0011010010101"  => dbus <= X"04C2EC8B";
				when "0011010010110"  => dbus <= X"97CE80C1";
				when "0011010010111"  => dbus <= X"D60397D6";
				when "0011010011000"  => dbus <= X"F0EF8267";
				when "0011010011001"  => dbus <= X"2783BF0F";
				when "0011010011010"  => dbus <= X"E0E300C0";
				when "0011010011011"  => dbus <= X"BBEDFEF4";
				when "0011010011100"  => dbus <= X"87936785";
				when "0011010011101"  => dbus <= X"08188207";
				when "0011010011110"  => dbus <= X"97BA79FD";
				when "0011010011111"  => dbus <= X"99BE4481";
				when "0011010100000"  => dbus <= X"04400A13";
				when "0011010100001"  => dbus <= X"2B376A85";
				when "0011010100010"  => dbus <= X"BFF14000";
				when "0011010100011"  => dbus <= X"034487B3";
				when "0011010100100"  => dbus <= X"048585A6";
				when "0011010100101"  => dbus <= X"EE4B0513";
				when "0011010100110"  => dbus <= X"80C104C2";
				when "0011010100111"  => dbus <= X"97D697CE";
				when "0011010101000"  => dbus <= X"8287D603";
				when "0011010101001"  => dbus <= X"BAEFF0EF";
				when "0011010101010"  => dbus <= X"00C02783";
				when "0011010101011"  => dbus <= X"FEF4E0E3";
				when "0011010101100"  => dbus <= X"6785B3C1";
				when "0011010101101"  => dbus <= X"82078793";
				when "0011010101110"  => dbus <= X"79FD0818";
				when "0011010101111"  => dbus <= X"448197BA";
				when "0011010110000"  => dbus <= X"0A1399BE";
				when "0011010110001"  => dbus <= X"6A850440";
				when "0011010110010"  => dbus <= X"40002B37";
				when "0011010110011"  => dbus <= X"87B3BFF1";
				when "0011010110100"  => dbus <= X"85A60344";
				when "0011010110101"  => dbus <= X"05130485";
				when "0011010110110"  => dbus <= X"04C2F00B";
				when "0011010110111"  => dbus <= X"97CE80C1";
				when "0011010111000"  => dbus <= X"D60397D6";
				when "0011010111001"  => dbus <= X"F0EF82A7";
				when "0011010111010"  => dbus <= X"2783B6CF";
				when "0011010111011"  => dbus <= X"E0E300C0";
				when "0011010111100"  => dbus <= X"B359FEF4";
				when "0011010111101"  => dbus <= X"87936785";
				when "0011010111110"  => dbus <= X"08188207";
				when "0011010111111"  => dbus <= X"97BA79FD";
				when "0011011000000"  => dbus <= X"99BE4481";
				when "0011011000001"  => dbus <= X"04400A13";
				when "0011011000010"  => dbus <= X"2B376A85";
				when "0011011000011"  => dbus <= X"BFF14000";
				when "0011011000100"  => dbus <= X"034487B3";
				when "0011011000101"  => dbus <= X"048585A6";
				when "0011011000110"  => dbus <= X"F1CB0513";
				when "0011011000111"  => dbus <= X"80C104C2";
				when "0011011001000"  => dbus <= X"97D697CE";
				when "0011011001001"  => dbus <= X"8247D603";
				when "0011011001010"  => dbus <= X"B2AFF0EF";
				when "0011011001011"  => dbus <= X"5763B39D";
				when "0011011001100"  => dbus <= X"25370080";
				when "0011011001101"  => dbus <= X"05134000";
				when "0011011001110"  => dbus <= X"B3B5F845";
				when "0011011001111"  => dbus <= X"40002537";
				when "0011011010000"  => dbus <= X"F9850513";
				when "0011011010001"  => dbus <= X"0000B38D";
				when "0011011010010"  => dbus <= X"3340D4B0";
				when "0011011010011"  => dbus <= X"E7146A79";
				when "0011011010100"  => dbus <= X"0000E3C1";
				when "0011011010101"  => dbus <= X"1199BE52";
				when "0011011010110"  => dbus <= X"1FD75608";
				when "0011011010111"  => dbus <= X"00000747";
				when "0011011011000"  => dbus <= X"39BF5E47";
				when "0011011011001"  => dbus <= X"8E3AE5A4";
				when "0011011011010"  => dbus <= X"00008D84";
				when "0011011011011"  => dbus <= X"40000970";
				when "0011011011100"  => dbus <= X"40000970";
				when "0011011011101"  => dbus <= X"40000976";
				when "0011011011110"  => dbus <= X"40000976";
				when "0011011011111"  => dbus <= X"4000097A";
				when "0011011100000"  => dbus <= X"40000A20";
				when "0011011100001"  => dbus <= X"400009FA";
				when "0011011100010"  => dbus <= X"40000A52";
				when "0011011100011"  => dbus <= X"40000ABE";
				when "0011011100100"  => dbus <= X"40000A78";
				when "0011011100101"  => dbus <= X"40000A98";
				when "0011011100110"  => dbus <= X"40000AD2";
				when "0011011100111"  => dbus <= X"40000AE8";
				when "0011011101000"  => dbus <= X"400020E0";
				when "0011011101001"  => dbus <= X"400020E8";
				when "0011011101010"  => dbus <= X"400020F0";
				when "0011011101011"  => dbus <= X"400020F8";
				when "0011011101100"  => dbus <= X"400020B0";
				when "0011011101101"  => dbus <= X"400020BC";
				when "0011011101110"  => dbus <= X"400020C8";
				when "0011011101111"  => dbus <= X"400020D4";
				when "0011011110000"  => dbus <= X"40002080";
				when "0011011110001"  => dbus <= X"4000208C";
				when "0011011110010"  => dbus <= X"40002098";
				when "0011011110011"  => dbus <= X"400020A4";
				when "0011011110100"  => dbus <= X"40002050";
				when "0011011110101"  => dbus <= X"4000205C";
				when "0011011110110"  => dbus <= X"40002068";
				when "0011011110111"  => dbus <= X"40002074";
				when "0011011111000"  => dbus <= X"40000C0A";
				when "0011011111001"  => dbus <= X"40000C10";
				when "0011011111010"  => dbus <= X"40000C16";
				when "0011011111011"  => dbus <= X"40000C1C";
				when "0011011111100"  => dbus <= X"40000C22";
				when "0011011111101"  => dbus <= X"70206B36";
				when "0011011111110"  => dbus <= X"6F667265";
				when "0011011111111"  => dbus <= X"6E616D72";
				when "0011100000000"  => dbus <= X"72206563";
				when "0011100000001"  => dbus <= X"70206E75";
				when "0011100000010"  => dbus <= X"6D617261";
				when "0011100000011"  => dbus <= X"72657465";
				when "0011100000100"  => dbus <= X"6F662073";
				when "0011100000101"  => dbus <= X"6F632072";
				when "0011100000110"  => dbus <= X"616D6572";
				when "0011100000111"  => dbus <= X"0A2E6B72";
				when "0011100001000"  => dbus <= X"00000000";
				when "0011100001001"  => dbus <= X"76206B36";
				when "0011100001010"  => dbus <= X"64696C61";
				when "0011100001011"  => dbus <= X"6F697461";
				when "0011100001100"  => dbus <= X"7572206E";
				when "0011100001101"  => dbus <= X"6170206E";
				when "0011100001110"  => dbus <= X"656D6172";
				when "0011100001111"  => dbus <= X"73726574";
				when "0011100010000"  => dbus <= X"726F6620";
				when "0011100010001"  => dbus <= X"726F6320";
				when "0011100010010"  => dbus <= X"72616D65";
				when "0011100010011"  => dbus <= X"000A2E6B";
				when "0011100010100"  => dbus <= X"666F7250";
				when "0011100010101"  => dbus <= X"20656C69";
				when "0011100010110"  => dbus <= X"656E6567";
				when "0011100010111"  => dbus <= X"69746172";
				when "0011100011000"  => dbus <= X"72206E6F";
				when "0011100011001"  => dbus <= X"70206E75";
				when "0011100011010"  => dbus <= X"6D617261";
				when "0011100011011"  => dbus <= X"72657465";
				when "0011100011100"  => dbus <= X"6F662073";
				when "0011100011101"  => dbus <= X"6F632072";
				when "0011100011110"  => dbus <= X"616D6572";
				when "0011100011111"  => dbus <= X"0A2E6B72";
				when "0011100100000"  => dbus <= X"00000000";
				when "0011100100001"  => dbus <= X"70204B32";
				when "0011100100010"  => dbus <= X"6F667265";
				when "0011100100011"  => dbus <= X"6E616D72";
				when "0011100100100"  => dbus <= X"72206563";
				when "0011100100101"  => dbus <= X"70206E75";
				when "0011100100110"  => dbus <= X"6D617261";
				when "0011100100111"  => dbus <= X"72657465";
				when "0011100101000"  => dbus <= X"6F662073";
				when "0011100101001"  => dbus <= X"6F632072";
				when "0011100101010"  => dbus <= X"616D6572";
				when "0011100101011"  => dbus <= X"0A2E6B72";
				when "0011100101100"  => dbus <= X"00000000";
				when "0011100101101"  => dbus <= X"76204B32";
				when "0011100101110"  => dbus <= X"64696C61";
				when "0011100101111"  => dbus <= X"6F697461";
				when "0011100110000"  => dbus <= X"7572206E";
				when "0011100110001"  => dbus <= X"6170206E";
				when "0011100110010"  => dbus <= X"656D6172";
				when "0011100110011"  => dbus <= X"73726574";
				when "0011100110100"  => dbus <= X"726F6620";
				when "0011100110101"  => dbus <= X"726F6320";
				when "0011100110110"  => dbus <= X"72616D65";
				when "0011100110111"  => dbus <= X"000A2E6B";
				when "0011100111000"  => dbus <= X"5D75255B";
				when "0011100111001"  => dbus <= X"4F525245";
				when "0011100111010"  => dbus <= X"6C202152";
				when "0011100111011"  => dbus <= X"20747369";
				when "0011100111100"  => dbus <= X"20637263";
				when "0011100111101"  => dbus <= X"30257830";
				when "0011100111110"  => dbus <= X"2D207834";
				when "0011100111111"  => dbus <= X"6F687320";
				when "0011101000000"  => dbus <= X"20646C75";
				when "0011101000001"  => dbus <= X"30206562";
				when "0011101000010"  => dbus <= X"34302578";
				when "0011101000011"  => dbus <= X"00000A78";
				when "0011101000100"  => dbus <= X"5D75255B";
				when "0011101000101"  => dbus <= X"4F525245";
				when "0011101000110"  => dbus <= X"6D202152";
				when "0011101000111"  => dbus <= X"69727461";
				when "0011101001000"  => dbus <= X"72632078";
				when "0011101001001"  => dbus <= X"78302063";
				when "0011101001010"  => dbus <= X"78343025";
				when "0011101001011"  => dbus <= X"73202D20";
				when "0011101001100"  => dbus <= X"6C756F68";
				when "0011101001101"  => dbus <= X"65622064";
				when "0011101001110"  => dbus <= X"25783020";
				when "0011101001111"  => dbus <= X"0A783430";
				when "0011101010000"  => dbus <= X"00000000";
				when "0011101010001"  => dbus <= X"5D75255B";
				when "0011101010010"  => dbus <= X"4F525245";
				when "0011101010011"  => dbus <= X"73202152";
				when "0011101010100"  => dbus <= X"65746174";
				when "0011101010101"  => dbus <= X"63726320";
				when "0011101010110"  => dbus <= X"25783020";
				when "0011101010111"  => dbus <= X"20783430";
				when "0011101011000"  => dbus <= X"6873202D";
				when "0011101011001"  => dbus <= X"646C756F";
				when "0011101011010"  => dbus <= X"20656220";
				when "0011101011011"  => dbus <= X"30257830";
				when "0011101011100"  => dbus <= X"000A7834";
				when "0011101011101"  => dbus <= X"65726F43";
				when "0011101011110"  => dbus <= X"6B72614D";
				when "0011101011111"  => dbus <= X"7A695320";
				when "0011101100000"  => dbus <= X"20202065";
				when "0011101100001"  => dbus <= X"25203A20";
				when "0011101100010"  => dbus <= X"000A756C";
				when "0011101100011"  => dbus <= X"61746F54";
				when "0011101100100"  => dbus <= X"6974206C";
				when "0011101100101"  => dbus <= X"20736B63";
				when "0011101100110"  => dbus <= X"20202020";
				when "0011101100111"  => dbus <= X"25203A20";
				when "0011101101000"  => dbus <= X"000A756C";
				when "0011101101001"  => dbus <= X"61746F54";
				when "0011101101010"  => dbus <= X"6974206C";
				when "0011101101011"  => dbus <= X"2820656D";
				when "0011101101100"  => dbus <= X"73636573";
				when "0011101101101"  => dbus <= X"25203A29";
				when "0011101101110"  => dbus <= X"00000A64";
				when "0011101101111"  => dbus <= X"72657449";
				when "0011101110000"  => dbus <= X"6F697461";
				when "0011101110001"  => dbus <= X"532F736E";
				when "0011101110010"  => dbus <= X"20206365";
				when "0011101110011"  => dbus <= X"25203A20";
				when "0011101110100"  => dbus <= X"00000A64";
				when "0011101110101"  => dbus <= X"4F525245";
				when "0011101110110"  => dbus <= X"4D202152";
				when "0011101110111"  => dbus <= X"20747375";
				when "0011101111000"  => dbus <= X"63657865";
				when "0011101111001"  => dbus <= X"20657475";
				when "0011101111010"  => dbus <= X"20726F66";
				when "0011101111011"  => dbus <= X"6C207461";
				when "0011101111100"  => dbus <= X"74736165";
				when "0011101111101"  => dbus <= X"20303120";
				when "0011101111110"  => dbus <= X"73636573";
				when "0011101111111"  => dbus <= X"726F6620";
				when "0011110000000"  => dbus <= X"76206120";
				when "0011110000001"  => dbus <= X"64696C61";
				when "0011110000010"  => dbus <= X"73657220";
				when "0011110000011"  => dbus <= X"21746C75";
				when "0011110000100"  => dbus <= X"0000000A";
				when "0011110000101"  => dbus <= X"72657449";
				when "0011110000110"  => dbus <= X"6F697461";
				when "0011110000111"  => dbus <= X"2020736E";
				when "0011110001000"  => dbus <= X"20202020";
				when "0011110001001"  => dbus <= X"25203A20";
				when "0011110001010"  => dbus <= X"000A756C";
				when "0011110001011"  => dbus <= X"38434347";
				when "0011110001100"  => dbus <= X"302E322E";
				when "0011110001101"  => dbus <= X"00000000";
				when "0011110001110"  => dbus <= X"706D6F43";
				when "0011110001111"  => dbus <= X"72656C69";
				when "0011110010000"  => dbus <= X"72657620";
				when "0011110010001"  => dbus <= X"6E6F6973";
				when "0011110010010"  => dbus <= X"25203A20";
				when "0011110010011"  => dbus <= X"00000A73";
				when "0011110010100"  => dbus <= X"20444D2D";
				when "0011110010101"  => dbus <= X"20734F2D";
				when "0011110010110"  => dbus <= X"62616D2D";
				when "0011110010111"  => dbus <= X"6C693D69";
				when "0011110011000"  => dbus <= X"20323370";
				when "0011110011001"  => dbus <= X"72616D2D";
				when "0011110011010"  => dbus <= X"723D6863";
				when "0011110011011"  => dbus <= X"69323376";
				when "0011110011100"  => dbus <= X"0000636D";
				when "0011110011101"  => dbus <= X"706D6F43";
				when "0011110011110"  => dbus <= X"72656C69";
				when "0011110011111"  => dbus <= X"616C6620";
				when "0011110100000"  => dbus <= X"20207367";
				when "0011110100001"  => dbus <= X"25203A20";
				when "0011110100010"  => dbus <= X"00000A73";
				when "0011110100011"  => dbus <= X"43415453";
				when "0011110100100"  => dbus <= X"0000004B";
				when "0011110100101"  => dbus <= X"6F6D654D";
				when "0011110100110"  => dbus <= X"6C207972";
				when "0011110100111"  => dbus <= X"7461636F";
				when "0011110101000"  => dbus <= X"206E6F69";
				when "0011110101001"  => dbus <= X"25203A20";
				when "0011110101010"  => dbus <= X"00000A73";
				when "0011110101011"  => dbus <= X"64656573";
				when "0011110101100"  => dbus <= X"20637263";
				when "0011110101101"  => dbus <= X"20202020";
				when "0011110101110"  => dbus <= X"20202020";
				when "0011110101111"  => dbus <= X"30203A20";
				when "0011110110000"  => dbus <= X"34302578";
				when "0011110110001"  => dbus <= X"00000A78";
				when "0011110110010"  => dbus <= X"5D64255B";
				when "0011110110011"  => dbus <= X"6C637263";
				when "0011110110100"  => dbus <= X"20747369";
				when "0011110110101"  => dbus <= X"20202020";
				when "0011110110110"  => dbus <= X"203A2020";
				when "0011110110111"  => dbus <= X"30257830";
				when "0011110111000"  => dbus <= X"000A7834";
				when "0011110111001"  => dbus <= X"5D64255B";
				when "0011110111010"  => dbus <= X"6D637263";
				when "0011110111011"  => dbus <= X"69727461";
				when "0011110111100"  => dbus <= X"20202078";
				when "0011110111101"  => dbus <= X"203A2020";
				when "0011110111110"  => dbus <= X"30257830";
				when "0011110111111"  => dbus <= X"000A7834";
				when "0011111000000"  => dbus <= X"5D64255B";
				when "0011111000001"  => dbus <= X"73637263";
				when "0011111000010"  => dbus <= X"65746174";
				when "0011111000011"  => dbus <= X"20202020";
				when "0011111000100"  => dbus <= X"203A2020";
				when "0011111000101"  => dbus <= X"30257830";
				when "0011111000110"  => dbus <= X"000A7834";
				when "0011111000111"  => dbus <= X"5D64255B";
				when "0011111001000"  => dbus <= X"66637263";
				when "0011111001001"  => dbus <= X"6C616E69";
				when "0011111001010"  => dbus <= X"20202020";
				when "0011111001011"  => dbus <= X"203A2020";
				when "0011111001100"  => dbus <= X"30257830";
				when "0011111001101"  => dbus <= X"000A7834";
				when "0011111001110"  => dbus <= X"72726F43";
				when "0011111001111"  => dbus <= X"20746365";
				when "0011111010000"  => dbus <= X"7265706F";
				when "0011111010001"  => dbus <= X"6F697461";
				when "0011111010010"  => dbus <= X"6176206E";
				when "0011111010011"  => dbus <= X"6164696C";
				when "0011111010100"  => dbus <= X"2E646574";
				when "0011111010101"  => dbus <= X"65655320";
				when "0011111010110"  => dbus <= X"41455220";
				when "0011111010111"  => dbus <= X"2E454D44";
				when "0011111011000"  => dbus <= X"6620646D";
				when "0011111011001"  => dbus <= X"7220726F";
				when "0011111011010"  => dbus <= X"61206E75";
				when "0011111011011"  => dbus <= X"7220646E";
				when "0011111011100"  => dbus <= X"726F7065";
				when "0011111011101"  => dbus <= X"676E6974";
				when "0011111011110"  => dbus <= X"6C757220";
				when "0011111011111"  => dbus <= X"0A2E7365";
				when "0011111100000"  => dbus <= X"00000000";
				when "0011111100001"  => dbus <= X"6F727245";
				when "0011111100010"  => dbus <= X"64207372";
				when "0011111100011"  => dbus <= X"63657465";
				when "0011111100100"  => dbus <= X"0A646574";
				when "0011111100101"  => dbus <= X"00000000";
				when "0011111100110"  => dbus <= X"6E6E6143";
				when "0011111100111"  => dbus <= X"7620746F";
				when "0011111101000"  => dbus <= X"64696C61";
				when "0011111101001"  => dbus <= X"20657461";
				when "0011111101010"  => dbus <= X"7265706F";
				when "0011111101011"  => dbus <= X"6F697461";
				when "0011111101100"  => dbus <= X"6F66206E";
				when "0011111101101"  => dbus <= X"68742072";
				when "0011111101110"  => dbus <= X"20657365";
				when "0011111101111"  => dbus <= X"64656573";
				when "0011111110000"  => dbus <= X"6C617620";
				when "0011111110001"  => dbus <= X"2C736575";
				when "0011111110010"  => dbus <= X"656C7020";
				when "0011111110011"  => dbus <= X"20657361";
				when "0011111110100"  => dbus <= X"706D6F63";
				when "0011111110101"  => dbus <= X"20657261";
				when "0011111110110"  => dbus <= X"68746977";
				when "0011111110111"  => dbus <= X"73657220";
				when "0011111111000"  => dbus <= X"73746C75";
				when "0011111111001"  => dbus <= X"206E6F20";
				when "0011111111010"  => dbus <= X"6E6B2061";
				when "0011111111011"  => dbus <= X"206E776F";
				when "0011111111100"  => dbus <= X"74616C70";
				when "0011111111101"  => dbus <= X"6D726F66";
				when "0011111111110"  => dbus <= X"00000A2E";
				when "0011111111111"  => dbus <= X"74617453";
				when "0100000000000"  => dbus <= X"00006369";
				when "0100000000001"  => dbus <= X"70616548";
				when "0100000000010"  => dbus <= X"00000000";
				when "0100000000011"  => dbus <= X"63617453";
				when "0100000000100"  => dbus <= X"0000006B";
				when "0100000000101"  => dbus <= X"72617453";
				when "0100000000110"  => dbus <= X"69742074";
				when "0100000000111"  => dbus <= X"2520656D";
				when "0100000001000"  => dbus <= X"000A646C";
				when "0100000001001"  => dbus <= X"706F7473";
				when "0100000001010"  => dbus <= X"6D697420";
				when "0100000001011"  => dbus <= X"6C252065";
				when "0100000001100"  => dbus <= X"00000A64";
				when "0100000001101"  => dbus <= X"72617453";
				when "0100000001110"  => dbus <= X"676E6974";
				when "0100000001111"  => dbus <= X"524F4320";
				when "0100000010000"  => dbus <= X"52414D45";
				when "0100000010001"  => dbus <= X"2E31204B";
				when "0100000010010"  => dbus <= X"2E2E2E30";
				when "0100000010011"  => dbus <= X"0000000A";
				when "0100000010100"  => dbus <= X"332E3054";
				when "0100000010101"  => dbus <= X"46312D65";
				when "0100000010110"  => dbus <= X"00000000";
				when "0100000010111"  => dbus <= X"542E542D";
				when "0100000011000"  => dbus <= X"71542B2B";
				when "0100000011001"  => dbus <= X"00000000";
				when "0100000011010"  => dbus <= X"2E335431";
				when "0100000011011"  => dbus <= X"7A346534";
				when "0100000011100"  => dbus <= X"00000000";
				when "0100000011101"  => dbus <= X"302E3433";
				when "0100000011110"  => dbus <= X"5E542D65";
				when "0100000011111"  => dbus <= X"00000000";
				when "0100000100000"  => dbus <= X"30352E35";
				when "0100000100001"  => dbus <= X"332B6530";
				when "0100000100010"  => dbus <= X"00000000";
				when "0100000100011"  => dbus <= X"32312E2D";
				when "0100000100100"  => dbus <= X"322D6533";
				when "0100000100101"  => dbus <= X"00000000";
				when "0100000100110"  => dbus <= X"6537382D";
				when "0100000100111"  => dbus <= X"3233382B";
				when "0100000101000"  => dbus <= X"00000000";
				when "0100000101001"  => dbus <= X"362E302B";
				when "0100000101010"  => dbus <= X"32312D65";
				when "0100000101011"  => dbus <= X"00000000";
				when "0100000101100"  => dbus <= X"352E3533";
				when "0100000101101"  => dbus <= X"30303434";
				when "0100000101110"  => dbus <= X"00000000";
				when "0100000101111"  => dbus <= X"3332312E";
				when "0100000110000"  => dbus <= X"30303534";
				when "0100000110001"  => dbus <= X"00000000";
				when "0100000110010"  => dbus <= X"3031312D";
				when "0100000110011"  => dbus <= X"3030372E";
				when "0100000110100"  => dbus <= X"00000000";
				when "0100000110101"  => dbus <= X"362E302B";
				when "0100000110110"  => dbus <= X"30303434";
				when "0100000110111"  => dbus <= X"00000000";
				when "0100000111000"  => dbus <= X"32313035";
				when "0100000111001"  => dbus <= X"00000000";
				when "0100000111010"  => dbus <= X"34333231";
				when "0100000111011"  => dbus <= X"00000000";
				when "0100000111100"  => dbus <= X"3437382D";
				when "0100000111101"  => dbus <= X"00000000";
				when "0100000111110"  => dbus <= X"3232312B";
				when "0100000111111"  => dbus <= X"00000000";
				when "0100001000000"  => dbus <= X"33323130";
				when "0100001000001"  => dbus <= X"37363534";
				when "0100001000010"  => dbus <= X"62613938";
				when "0100001000011"  => dbus <= X"66656463";
				when "0100001000100"  => dbus <= X"6A696867";
				when "0100001000101"  => dbus <= X"6E6D6C6B";
				when "0100001000110"  => dbus <= X"7271706F";
				when "0100001000111"  => dbus <= X"76757473";
				when "0100001001000"  => dbus <= X"7A797877";
				when "0100001001001"  => dbus <= X"00000000";
				when "0100001001010"  => dbus <= X"33323130";
				when "0100001001011"  => dbus <= X"37363534";
				when "0100001001100"  => dbus <= X"42413938";
				when "0100001001101"  => dbus <= X"46454443";
				when "0100001001110"  => dbus <= X"4A494847";
				when "0100001001111"  => dbus <= X"4E4D4C4B";
				when "0100001010000"  => dbus <= X"5251504F";
				when "0100001010001"  => dbus <= X"56555453";
				when "0100001010010"  => dbus <= X"5A595857";
				when "0100001010011"  => dbus <= X"00000000";
				when "0100001010100"  => dbus <= X"4C554E3C";
				when "0100001010101"  => dbus <= X"00003E4C";
				when "0100001010110"  => dbus <= X"33323130";
				when "0100001010111"  => dbus <= X"37363534";
				when "0100001011000"  => dbus <= X"42413938";
				when "0100001011001"  => dbus <= X"46454443";
				when "0100001011010"  => dbus <= X"00000000";
				when "0100001011011"  => dbus <= X"40001FFC";
				when "0100001011100"  => dbus <= X"40002004";
				when "0100001011101"  => dbus <= X"4000200C";
				when "0100001011110"  => dbus <= X"00000001";
				when "0100001011111"  => dbus <= X"00000001";
				when "0100001100000"  => dbus <= X"00000066";
				when "0100001100001"  => dbus <= X"00000066";
				when others    => dbus <= "00000000000000000000000000000000";
				end case;
			end if;
		end if;
	end process;
end rtl;
