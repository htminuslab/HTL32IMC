-------------------------------------------------------------------------------
--  HTLROM32                                                                 --
--  Copyright (C) 2002-2025 HT-LAB                                           --
--                                                                           --
-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- Project       :                                                           --
-- Purpose       :                                                           --
-- Library       :                                                           --
--                                                                           --
-- Created       : bin2text -vhd version  0.5                                --
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.ALL;

entity bootloader is
	port(clk    : in  std_logic;
		 abus   : in  std_logic_vector(12 downto 0);
		 ena    : in std_logic;
		 dbus   : out std_logic_vector(31 downto 0));
end bootloader;

architecture rtl of bootloader is
begin

	process(clk)
		begin
		if rising_edge(clk) then
			if ena='1' then
			case abus is
				when "0000000000000"  => dbus <= X"0100006F";
				when "0000000000001"  => dbus <= X"00000013";
				when "0000000000010"  => dbus <= X"00000013";
				when "0000000000011"  => dbus <= X"00000013";
				when "0000000000100"  => dbus <= X"00008137";
				when "0000000000101"  => dbus <= X"B8010113";
				when "0000000000110"  => dbus <= X"00000517";
				when "0000000000111"  => dbus <= X"41050513";
				when "0000000001000"  => dbus <= X"00000593";
				when "0000000001001"  => dbus <= X"00000613";
				when "0000000001010"  => dbus <= X"00C5DC63";
				when "0000000001011"  => dbus <= X"00052683";
				when "0000000001100"  => dbus <= X"00D5A023";
				when "0000000001101"  => dbus <= X"00450513";
				when "0000000001110"  => dbus <= X"00458593";
				when "0000000001111"  => dbus <= X"FEC5C8E3";
				when "0000000010000"  => dbus <= X"00000513";
				when "0000000010001"  => dbus <= X"00800593";
				when "0000000010010"  => dbus <= X"00B55863";
				when "0000000010011"  => dbus <= X"00052023";
				when "0000000010100"  => dbus <= X"00450513";
				when "0000000010101"  => dbus <= X"FEB54CE3";
				when "0000000010110"  => dbus <= X"330000EF";
				when "0000000010111"  => dbus <= X"00100073";
				when "0000000011000"  => dbus <= X"00000793";
				when "0000000011001"  => dbus <= X"00C79463";
				when "0000000011010"  => dbus <= X"00008067";
				when "0000000011011"  => dbus <= X"00F58733";
				when "0000000011100"  => dbus <= X"00074683";
				when "0000000011101"  => dbus <= X"00F50733";
				when "0000000011110"  => dbus <= X"00178793";
				when "0000000011111"  => dbus <= X"00D70023";
				when "0000000100000"  => dbus <= X"FE5FF06F";
				when "0000000100001"  => dbus <= X"800007B7";
				when "0000000100010"  => dbus <= X"08A78023";
				when "0000000100011"  => dbus <= X"00008067";
				when "0000000100100"  => dbus <= X"80000737";
				when "0000000100101"  => dbus <= X"00054783";
				when "0000000100110"  => dbus <= X"00079463";
				when "0000000100111"  => dbus <= X"00008067";
				when "0000000101000"  => dbus <= X"00150513";
				when "0000000101001"  => dbus <= X"08F70023";
				when "0000000101010"  => dbus <= X"FEDFF06F";
				when "0000000101011"  => dbus <= X"FF010113";
				when "0000000101100"  => dbus <= X"00410793";
				when "0000000101101"  => dbus <= X"00078693";
				when "0000000101110"  => dbus <= X"00A00713";
				when "0000000101111"  => dbus <= X"02051663";
				when "0000000110000"  => dbus <= X"02D78463";
				when "0000000110001"  => dbus <= X"80000637";
				when "0000000110010"  => dbus <= X"FFF78793";
				when "0000000110011"  => dbus <= X"0007C703";
				when "0000000110100"  => dbus <= X"03070713";
				when "0000000110101"  => dbus <= X"0FF77713";
				when "0000000110110"  => dbus <= X"08E60023";
				when "0000000110111"  => dbus <= X"FED796E3";
				when "0000000111000"  => dbus <= X"01010113";
				when "0000000111001"  => dbus <= X"00008067";
				when "0000000111010"  => dbus <= X"02E57633";
				when "0000000111011"  => dbus <= X"00178793";
				when "0000000111100"  => dbus <= X"FEC78FA3";
				when "0000000111101"  => dbus <= X"02E55533";
				when "0000000111110"  => dbus <= X"FC5FF06F";
				when "0000000111111"  => dbus <= X"FFF58593";
				when "0000001000000"  => dbus <= X"40000737";
				when "0000001000001"  => dbus <= X"00259593";
				when "0000001000010"  => dbus <= X"3E070713";
				when "0000001000011"  => dbus <= X"800006B7";
				when "0000001000100"  => dbus <= X"0005D463";
				when "0000001000101"  => dbus <= X"00008067";
				when "0000001000110"  => dbus <= X"00B557B3";
				when "0000001000111"  => dbus <= X"00F7F793";
				when "0000001001000"  => dbus <= X"00E787B3";
				when "0000001001001"  => dbus <= X"0007C783";
				when "0000001001010"  => dbus <= X"FFC58593";
				when "0000001001011"  => dbus <= X"08F68023";
				when "0000001001100"  => dbus <= X"FE1FF06F";
				when "0000001001101"  => dbus <= X"80000737";
				when "0000001001110"  => dbus <= X"00C72783";
				when "0000001001111"  => dbus <= X"0017F793";
				when "0000001010000"  => dbus <= X"FE078CE3";
				when "0000001010001"  => dbus <= X"00A72223";
				when "0000001010010"  => dbus <= X"00008067";
				when "0000001010011"  => dbus <= X"80000737";
				when "0000001010100"  => dbus <= X"00C72783";
				when "0000001010101"  => dbus <= X"0027F793";
				when "0000001010110"  => dbus <= X"FE078CE3";
				when "0000001010111"  => dbus <= X"00072503";
				when "0000001011000"  => dbus <= X"0FF57513";
				when "0000001011001"  => dbus <= X"00008067";
				when "0000001011010"  => dbus <= X"80000737";
				when "0000001011011"  => dbus <= X"01C72783";
				when "0000001011100"  => dbus <= X"0017F793";
				when "0000001011101"  => dbus <= X"FE078CE3";
				when "0000001011110"  => dbus <= X"00A72A23";
				when "0000001011111"  => dbus <= X"00008067";
				when "0000001100000"  => dbus <= X"80000737";
				when "0000001100001"  => dbus <= X"01C72783";
				when "0000001100010"  => dbus <= X"0027F793";
				when "0000001100011"  => dbus <= X"FE078CE3";
				when "0000001100100"  => dbus <= X"01072503";
				when "0000001100101"  => dbus <= X"0FF57513";
				when "0000001100110"  => dbus <= X"00008067";
				when "0000001100111"  => dbus <= X"FF010113";
				when "0000001101000"  => dbus <= X"00812423";
				when "0000001101001"  => dbus <= X"00112623";
				when "0000001101010"  => dbus <= X"00050413";
				when "0000001101011"  => dbus <= X"00044503";
				when "0000001101100"  => dbus <= X"00051A63";
				when "0000001101101"  => dbus <= X"00C12083";
				when "0000001101110"  => dbus <= X"00812403";
				when "0000001101111"  => dbus <= X"01010113";
				when "0000001110000"  => dbus <= X"00008067";
				when "0000001110001"  => dbus <= X"00140413";
				when "0000001110010"  => dbus <= X"F6DFF0EF";
				when "0000001110011"  => dbus <= X"FE1FF06F";
				when "0000001110100"  => dbus <= X"FF010113";
				when "0000001110101"  => dbus <= X"00812423";
				when "0000001110110"  => dbus <= X"00112623";
				when "0000001110111"  => dbus <= X"00050413";
				when "0000001111000"  => dbus <= X"00044503";
				when "0000001111001"  => dbus <= X"00051A63";
				when "0000001111010"  => dbus <= X"00C12083";
				when "0000001111011"  => dbus <= X"00812403";
				when "0000001111100"  => dbus <= X"01010113";
				when "0000001111101"  => dbus <= X"00008067";
				when "0000001111110"  => dbus <= X"00140413";
				when "0000001111111"  => dbus <= X"F6DFF0EF";
				when "0000010000000"  => dbus <= X"FE1FF06F";
				when "0000010000001"  => dbus <= X"C81027F3";
				when "0000010000010"  => dbus <= X"C0102573";
				when "0000010000011"  => dbus <= X"C81025F3";
				when "0000010000100"  => dbus <= X"FEF59AE3";
				when "0000010000101"  => dbus <= X"00008067";
				when "0000010000110"  => dbus <= X"FF010113";
				when "0000010000111"  => dbus <= X"00812423";
				when "0000010001000"  => dbus <= X"00912223";
				when "0000010001001"  => dbus <= X"00112623";
				when "0000010001010"  => dbus <= X"00050413";
				when "0000010001011"  => dbus <= X"00058493";
				when "0000010001100"  => dbus <= X"FD5FF0EF";
				when "0000010001101"  => dbus <= X"008507B3";
				when "0000010001110"  => dbus <= X"00A7B533";
				when "0000010001111"  => dbus <= X"009585B3";
				when "0000010010000"  => dbus <= X"00B50533";
				when "0000010010001"  => dbus <= X"FFF00713";
				when "0000010010010"  => dbus <= X"88371073";
				when "0000010010011"  => dbus <= X"80379073";
				when "0000010010100"  => dbus <= X"88351073";
				when "0000010010101"  => dbus <= X"00C12083";
				when "0000010010110"  => dbus <= X"00812403";
				when "0000010010111"  => dbus <= X"00412483";
				when "0000010011000"  => dbus <= X"01010113";
				when "0000010011001"  => dbus <= X"00008067";
				when "0000010011010"  => dbus <= X"FB010113";
				when "0000010011011"  => dbus <= X"04112623";
				when "0000010011100"  => dbus <= X"04512423";
				when "0000010011101"  => dbus <= X"04612223";
				when "0000010011110"  => dbus <= X"04712023";
				when "0000010011111"  => dbus <= X"02812E23";
				when "0000010100000"  => dbus <= X"02912C23";
				when "0000010100001"  => dbus <= X"02A12A23";
				when "0000010100010"  => dbus <= X"02B12823";
				when "0000010100011"  => dbus <= X"02C12623";
				when "0000010100100"  => dbus <= X"02D12423";
				when "0000010100101"  => dbus <= X"02E12223";
				when "0000010100110"  => dbus <= X"02F12023";
				when "0000010100111"  => dbus <= X"01012E23";
				when "0000010101000"  => dbus <= X"01112C23";
				when "0000010101001"  => dbus <= X"01C12A23";
				when "0000010101010"  => dbus <= X"01D12823";
				when "0000010101011"  => dbus <= X"01E12623";
				when "0000010101100"  => dbus <= X"01F12423";
				when "0000010101101"  => dbus <= X"34202473";
				when "0000010101110"  => dbus <= X"800007B7";
				when "0000010101111"  => dbus <= X"400004B7";
				when "0000010110000"  => dbus <= X"0AF41663";
				when "0000010110001"  => dbus <= X"00002503";
				when "0000010110010"  => dbus <= X"000017B7";
				when "0000010110011"  => dbus <= X"00402583";
				when "0000010110100"  => dbus <= X"77078793";
				when "0000010110101"  => dbus <= X"00F507B3";
				when "0000010110110"  => dbus <= X"00A7B733";
				when "0000010110111"  => dbus <= X"00F02023";
				when "0000010111000"  => dbus <= X"00B706B3";
				when "0000010111001"  => dbus <= X"00D02223";
				when "0000010111010"  => dbus <= X"00002503";
				when "0000010111011"  => dbus <= X"00402583";
				when "0000010111100"  => dbus <= X"F29FF0EF";
				when "0000010111101"  => dbus <= X"40000537";
				when "0000010111110"  => dbus <= X"3F450513";
				when "0000010111111"  => dbus <= X"D95FF0EF";
				when "0000011000000"  => dbus <= X"00002783";
				when "0000011000001"  => dbus <= X"00402803";
				when "0000011000010"  => dbus <= X"00800593";
				when "0000011000011"  => dbus <= X"00078513";
				when "0000011000100"  => dbus <= X"DEDFF0EF";
				when "0000011000101"  => dbus <= X"40048513";
				when "0000011000110"  => dbus <= X"D79FF0EF";
				when "0000011000111"  => dbus <= X"03C12403";
				when "0000011001000"  => dbus <= X"04C12083";
				when "0000011001001"  => dbus <= X"04812283";
				when "0000011001010"  => dbus <= X"04412303";
				when "0000011001011"  => dbus <= X"04012383";
				when "0000011001100"  => dbus <= X"03812483";
				when "0000011001101"  => dbus <= X"03412503";
				when "0000011001110"  => dbus <= X"03012583";
				when "0000011001111"  => dbus <= X"02C12603";
				when "0000011010000"  => dbus <= X"02812683";
				when "0000011010001"  => dbus <= X"02412703";
				when "0000011010010"  => dbus <= X"02012783";
				when "0000011010011"  => dbus <= X"01C12803";
				when "0000011010100"  => dbus <= X"01812883";
				when "0000011010101"  => dbus <= X"01412E03";
				when "0000011010110"  => dbus <= X"01012E83";
				when "0000011010111"  => dbus <= X"00C12F03";
				when "0000011011000"  => dbus <= X"00812F83";
				when "0000011011001"  => dbus <= X"05010113";
				when "0000011011010"  => dbus <= X"30200073";
				when "0000011011011"  => dbus <= X"40000537";
				when "0000011011100"  => dbus <= X"40450513";
				when "0000011011101"  => dbus <= X"D1DFF0EF";
				when "0000011011110"  => dbus <= X"00445513";
				when "0000011011111"  => dbus <= X"00357513";
				when "0000011100000"  => dbus <= X"D2DFF0EF";
				when "0000011100001"  => dbus <= X"F91FF06F";
				when "0000011100010"  => dbus <= X"40000537";
				when "0000011100011"  => dbus <= X"FF010113";
				when "0000011100100"  => dbus <= X"41850513";
				when "0000011100101"  => dbus <= X"00112623";
				when "0000011100110"  => dbus <= X"CF9FF0EF";
				when "0000011100111"  => dbus <= X"E69FF0EF";
				when "0000011101000"  => dbus <= X"000017B7";
				when "0000011101001"  => dbus <= X"77078793";
				when "0000011101010"  => dbus <= X"00F507B3";
				when "0000011101011"  => dbus <= X"00A7B733";
				when "0000011101100"  => dbus <= X"00B705B3";
				when "0000011101101"  => dbus <= X"00078513";
				when "0000011101110"  => dbus <= X"E61FF0EF";
				when "0000011101111"  => dbus <= X"400007B7";
				when "0000011110000"  => dbus <= X"26878793";
				when "0000011110001"  => dbus <= X"30579073";
				when "0000011110010"  => dbus <= X"08000793";
				when "0000011110011"  => dbus <= X"30479073";
				when "0000011110100"  => dbus <= X"00800793";
				when "0000011110101"  => dbus <= X"30079073";
				when "0000011110110"  => dbus <= X"10500073";
				when "0000011110111"  => dbus <= X"FFDFF06F";
				when "0000011111000"  => dbus <= X"33323130";
				when "0000011111001"  => dbus <= X"37363534";
				when "0000011111010"  => dbus <= X"42413938";
				when "0000011111011"  => dbus <= X"46454443";
				when "0000011111100"  => dbus <= X"00000000";
				when "0000011111101"  => dbus <= X"5152490A";
				when "0000011111110"  => dbus <= X"524D5420";
				when "0000011111111"  => dbus <= X"0000003D";
				when "0000100000000"  => dbus <= X"0000000A";
				when "0000100000001"  => dbus <= X"3E3E3E3E";
				when "0000100000010"  => dbus <= X"74784520";
				when "0000100000011"  => dbus <= X"616E7265";
				when "0000100000100"  => dbus <= X"5249206C";
				when "0000100000101"  => dbus <= X"00000051";
				when "0000100000110"  => dbus <= X"656D6954";
				when "0000100000111"  => dbus <= X"52492072";
				when "0000100001000"  => dbus <= X"65542051";
				when "0000100001001"  => dbus <= X"000A7473";
				when "0000100001010"  => dbus <= X"000A7473";
				when others    => dbus <= "00000000000000000000000000000000";
				end case;
			end if;
		end if;
	end process;
end rtl;
